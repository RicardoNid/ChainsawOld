// Generator : SpinalHDL v1.4.2    git head : 804c7bd7b7feaddcc1d25ecef6c208fd5f776f79
// Component : FIR
// Git hash  : faa40885e164272f61221e4440a1cea60f1bc866



module FIR (
  input      [26:0]   io_dataIn,
  output     [47:0]   io_dataOut,
  input               clk,
  input               reset
);
  wire       [47:0]   _zz_289;
  wire       [47:0]   _zz_290;
  wire       [47:0]   _zz_291;
  wire       [47:0]   _zz_292;
  wire       [47:0]   _zz_293;
  wire       [47:0]   _zz_294;
  wire       [47:0]   _zz_295;
  wire       [47:0]   _zz_296;
  wire       [47:0]   _zz_297;
  wire       [47:0]   _zz_298;
  wire       [47:0]   _zz_299;
  wire       [47:0]   _zz_300;
  wire       [47:0]   _zz_301;
  wire       [47:0]   _zz_302;
  wire       [47:0]   _zz_303;
  wire       [47:0]   _zz_304;
  wire       [47:0]   _zz_305;
  wire       [47:0]   _zz_306;
  wire       [47:0]   _zz_307;
  wire       [47:0]   _zz_308;
  wire       [47:0]   _zz_309;
  wire       [47:0]   _zz_310;
  wire       [47:0]   _zz_311;
  wire       [47:0]   _zz_312;
  wire       [47:0]   _zz_313;
  wire       [47:0]   _zz_314;
  wire       [47:0]   _zz_315;
  wire       [47:0]   _zz_316;
  wire       [47:0]   _zz_317;
  wire       [47:0]   _zz_318;
  wire       [47:0]   _zz_319;
  wire       [47:0]   _zz_320;
  wire       [47:0]   _zz_321;
  wire       [47:0]   _zz_322;
  wire       [47:0]   _zz_323;
  wire       [47:0]   _zz_324;
  wire       [47:0]   _zz_325;
  wire       [47:0]   _zz_326;
  wire       [47:0]   _zz_327;
  wire       [47:0]   _zz_328;
  wire       [47:0]   _zz_329;
  wire       [47:0]   _zz_330;
  wire       [47:0]   _zz_331;
  wire       [47:0]   _zz_332;
  wire       [47:0]   _zz_333;
  wire       [47:0]   _zz_334;
  wire       [47:0]   _zz_335;
  wire       [47:0]   _zz_336;
  wire       [47:0]   _zz_337;
  wire       [47:0]   _zz_338;
  wire       [47:0]   _zz_339;
  wire       [47:0]   _zz_340;
  wire       [47:0]   _zz_341;
  wire       [47:0]   _zz_342;
  wire       [47:0]   _zz_343;
  wire       [47:0]   _zz_344;
  wire       [47:0]   _zz_345;
  wire       [47:0]   _zz_346;
  wire       [47:0]   _zz_347;
  wire       [47:0]   _zz_348;
  wire       [47:0]   _zz_349;
  wire       [47:0]   _zz_350;
  wire       [47:0]   _zz_351;
  wire       [47:0]   _zz_352;
  wire       [47:0]   _zz_353;
  wire       [47:0]   _zz_354;
  wire       [47:0]   _zz_355;
  wire       [47:0]   _zz_356;
  wire       [47:0]   _zz_357;
  wire       [47:0]   _zz_358;
  wire       [47:0]   _zz_359;
  wire       [17:0]   weightWires_0;
  wire       [17:0]   weightWires_1;
  wire       [17:0]   weightWires_2;
  wire       [17:0]   weightWires_3;
  wire       [17:0]   weightWires_4;
  wire       [17:0]   weightWires_5;
  wire       [17:0]   weightWires_6;
  wire       [17:0]   weightWires_7;
  wire       [17:0]   weightWires_8;
  wire       [17:0]   weightWires_9;
  wire       [17:0]   weightWires_10;
  wire       [17:0]   weightWires_11;
  wire       [17:0]   weightWires_12;
  wire       [17:0]   weightWires_13;
  wire       [17:0]   weightWires_14;
  wire       [17:0]   weightWires_15;
  wire       [17:0]   weightWires_16;
  wire       [17:0]   weightWires_17;
  wire       [17:0]   weightWires_18;
  wire       [17:0]   weightWires_19;
  wire       [17:0]   weightWires_20;
  wire       [17:0]   weightWires_21;
  wire       [17:0]   weightWires_22;
  wire       [17:0]   weightWires_23;
  wire       [17:0]   weightWires_24;
  wire       [17:0]   weightWires_25;
  wire       [17:0]   weightWires_26;
  wire       [17:0]   weightWires_27;
  wire       [17:0]   weightWires_28;
  wire       [17:0]   weightWires_29;
  wire       [17:0]   weightWires_30;
  wire       [17:0]   weightWires_31;
  wire       [17:0]   weightWires_32;
  wire       [17:0]   weightWires_33;
  wire       [17:0]   weightWires_34;
  wire       [17:0]   weightWires_35;
  wire       [17:0]   weightWires_36;
  wire       [17:0]   weightWires_37;
  wire       [17:0]   weightWires_38;
  wire       [17:0]   weightWires_39;
  wire       [17:0]   weightWires_40;
  wire       [17:0]   weightWires_41;
  wire       [17:0]   weightWires_42;
  wire       [17:0]   weightWires_43;
  wire       [17:0]   weightWires_44;
  wire       [17:0]   weightWires_45;
  wire       [17:0]   weightWires_46;
  wire       [17:0]   weightWires_47;
  wire       [17:0]   weightWires_48;
  wire       [17:0]   weightWires_49;
  wire       [17:0]   weightWires_50;
  wire       [17:0]   weightWires_51;
  wire       [17:0]   weightWires_52;
  wire       [17:0]   weightWires_53;
  wire       [17:0]   weightWires_54;
  wire       [17:0]   weightWires_55;
  wire       [17:0]   weightWires_56;
  wire       [17:0]   weightWires_57;
  wire       [17:0]   weightWires_58;
  wire       [17:0]   weightWires_59;
  wire       [17:0]   weightWires_60;
  wire       [17:0]   weightWires_61;
  wire       [17:0]   weightWires_62;
  wire       [17:0]   weightWires_63;
  wire       [17:0]   weightWires_64;
  wire       [17:0]   weightWires_65;
  wire       [17:0]   weightWires_66;
  wire       [17:0]   weightWires_67;
  wire       [17:0]   weightWires_68;
  wire       [17:0]   weightWires_69;
  wire       [17:0]   weightWires_70;
  wire       [17:0]   weightWires_71;
  wire       [26:0]   inputZERO;
  reg        [26:0]   io_dataIn_regNext;
  reg        [26:0]   _zz_1;
  reg        [26:0]   _zz_2;
  reg        [26:0]   _zz_3;
  reg        [26:0]   _zz_4;
  reg        [26:0]   _zz_5;
  reg        [26:0]   _zz_6;
  reg        [26:0]   _zz_7;
  reg        [26:0]   _zz_8;
  reg        [26:0]   _zz_9;
  reg        [26:0]   _zz_10;
  reg        [26:0]   _zz_11;
  reg        [26:0]   _zz_12;
  reg        [26:0]   _zz_13;
  reg        [26:0]   _zz_14;
  reg        [26:0]   _zz_15;
  reg        [26:0]   _zz_16;
  reg        [26:0]   _zz_17;
  reg        [26:0]   _zz_18;
  reg        [26:0]   _zz_19;
  reg        [26:0]   _zz_20;
  reg        [26:0]   _zz_21;
  reg        [26:0]   _zz_22;
  reg        [26:0]   _zz_23;
  reg        [26:0]   _zz_24;
  reg        [26:0]   _zz_25;
  reg        [26:0]   _zz_26;
  reg        [26:0]   _zz_27;
  reg        [26:0]   _zz_28;
  reg        [26:0]   _zz_29;
  reg        [26:0]   _zz_30;
  reg        [26:0]   _zz_31;
  reg        [26:0]   _zz_32;
  reg        [26:0]   _zz_33;
  reg        [26:0]   _zz_34;
  reg        [26:0]   _zz_35;
  reg        [26:0]   _zz_36;
  reg        [26:0]   _zz_37;
  reg        [26:0]   _zz_38;
  reg        [26:0]   _zz_39;
  reg        [26:0]   _zz_40;
  reg        [26:0]   _zz_41;
  reg        [26:0]   _zz_42;
  reg        [26:0]   _zz_43;
  reg        [26:0]   _zz_44;
  reg        [26:0]   _zz_45;
  reg        [26:0]   _zz_46;
  reg        [26:0]   _zz_47;
  reg        [26:0]   _zz_48;
  reg        [26:0]   _zz_49;
  reg        [26:0]   _zz_50;
  reg        [26:0]   _zz_51;
  reg        [26:0]   _zz_52;
  reg        [26:0]   _zz_53;
  reg        [26:0]   _zz_54;
  reg        [26:0]   _zz_55;
  reg        [26:0]   _zz_56;
  reg        [26:0]   _zz_57;
  reg        [26:0]   _zz_58;
  reg        [26:0]   _zz_59;
  reg        [26:0]   _zz_60;
  reg        [26:0]   _zz_61;
  reg        [26:0]   _zz_62;
  reg        [26:0]   _zz_63;
  reg        [26:0]   _zz_64;
  reg        [26:0]   _zz_65;
  reg        [26:0]   _zz_66;
  reg        [26:0]   _zz_67;
  reg        [26:0]   _zz_68;
  reg        [26:0]   _zz_69;
  reg        [26:0]   _zz_70;
  reg        [26:0]   _zz_71;
  reg        [26:0]   _zz_72;
  reg        [26:0]   _zz_73;
  reg        [26:0]   _zz_74;
  reg        [26:0]   _zz_75;
  reg        [26:0]   _zz_76;
  reg        [26:0]   _zz_77;
  reg        [26:0]   _zz_78;
  reg        [26:0]   _zz_79;
  reg        [26:0]   _zz_80;
  reg        [26:0]   _zz_81;
  reg        [26:0]   _zz_82;
  reg        [26:0]   _zz_83;
  reg        [26:0]   _zz_84;
  reg        [26:0]   _zz_85;
  reg        [26:0]   _zz_86;
  reg        [26:0]   _zz_87;
  reg        [26:0]   _zz_88;
  reg        [26:0]   _zz_89;
  reg        [26:0]   _zz_90;
  reg        [26:0]   _zz_91;
  reg        [26:0]   _zz_92;
  reg        [26:0]   _zz_93;
  reg        [26:0]   _zz_94;
  reg        [26:0]   _zz_95;
  reg        [26:0]   _zz_96;
  reg        [26:0]   _zz_97;
  reg        [26:0]   _zz_98;
  reg        [26:0]   _zz_99;
  reg        [26:0]   _zz_100;
  reg        [26:0]   _zz_101;
  reg        [26:0]   _zz_102;
  reg        [26:0]   _zz_103;
  reg        [26:0]   _zz_104;
  reg        [26:0]   _zz_105;
  reg        [26:0]   _zz_106;
  reg        [26:0]   _zz_107;
  reg        [26:0]   _zz_108;
  reg        [26:0]   _zz_109;
  reg        [26:0]   _zz_110;
  reg        [26:0]   _zz_111;
  reg        [26:0]   _zz_112;
  reg        [26:0]   _zz_113;
  reg        [26:0]   _zz_114;
  reg        [26:0]   _zz_115;
  reg        [26:0]   _zz_116;
  reg        [26:0]   _zz_117;
  reg        [26:0]   _zz_118;
  reg        [26:0]   _zz_119;
  reg        [26:0]   _zz_120;
  reg        [26:0]   _zz_121;
  reg        [26:0]   _zz_122;
  reg        [26:0]   _zz_123;
  reg        [26:0]   _zz_124;
  reg        [26:0]   _zz_125;
  reg        [26:0]   _zz_126;
  reg        [26:0]   _zz_127;
  reg        [26:0]   _zz_128;
  reg        [26:0]   _zz_129;
  reg        [26:0]   _zz_130;
  reg        [26:0]   _zz_131;
  reg        [26:0]   _zz_132;
  reg        [26:0]   _zz_133;
  reg        [26:0]   _zz_134;
  reg        [26:0]   _zz_135;
  reg        [26:0]   _zz_136;
  reg        [26:0]   _zz_137;
  reg        [26:0]   _zz_138;
  reg        [26:0]   _zz_139;
  reg        [26:0]   _zz_140;
  reg        [26:0]   _zz_141;
  reg        [26:0]   _zz_142;
  reg        [26:0]   _zz_143;
  reg        [44:0]   _zz_144;
  reg        [44:0]   _zz_145;
  reg        [44:0]   _zz_146;
  reg        [44:0]   _zz_147;
  reg        [44:0]   _zz_148;
  reg        [44:0]   _zz_149;
  reg        [44:0]   _zz_150;
  reg        [44:0]   _zz_151;
  reg        [44:0]   _zz_152;
  reg        [44:0]   _zz_153;
  reg        [44:0]   _zz_154;
  reg        [44:0]   _zz_155;
  reg        [44:0]   _zz_156;
  reg        [44:0]   _zz_157;
  reg        [44:0]   _zz_158;
  reg        [44:0]   _zz_159;
  reg        [44:0]   _zz_160;
  reg        [44:0]   _zz_161;
  reg        [44:0]   _zz_162;
  reg        [44:0]   _zz_163;
  reg        [44:0]   _zz_164;
  reg        [44:0]   _zz_165;
  reg        [44:0]   _zz_166;
  reg        [44:0]   _zz_167;
  reg        [44:0]   _zz_168;
  reg        [44:0]   _zz_169;
  reg        [44:0]   _zz_170;
  reg        [44:0]   _zz_171;
  reg        [44:0]   _zz_172;
  reg        [44:0]   _zz_173;
  reg        [44:0]   _zz_174;
  reg        [44:0]   _zz_175;
  reg        [44:0]   _zz_176;
  reg        [44:0]   _zz_177;
  reg        [44:0]   _zz_178;
  reg        [44:0]   _zz_179;
  reg        [44:0]   _zz_180;
  reg        [44:0]   _zz_181;
  reg        [44:0]   _zz_182;
  reg        [44:0]   _zz_183;
  reg        [44:0]   _zz_184;
  reg        [44:0]   _zz_185;
  reg        [44:0]   _zz_186;
  reg        [44:0]   _zz_187;
  reg        [44:0]   _zz_188;
  reg        [44:0]   _zz_189;
  reg        [44:0]   _zz_190;
  reg        [44:0]   _zz_191;
  reg        [44:0]   _zz_192;
  reg        [44:0]   _zz_193;
  reg        [44:0]   _zz_194;
  reg        [44:0]   _zz_195;
  reg        [44:0]   _zz_196;
  reg        [44:0]   _zz_197;
  reg        [44:0]   _zz_198;
  reg        [44:0]   _zz_199;
  reg        [44:0]   _zz_200;
  reg        [44:0]   _zz_201;
  reg        [44:0]   _zz_202;
  reg        [44:0]   _zz_203;
  reg        [44:0]   _zz_204;
  reg        [44:0]   _zz_205;
  reg        [44:0]   _zz_206;
  reg        [44:0]   _zz_207;
  reg        [44:0]   _zz_208;
  reg        [44:0]   _zz_209;
  reg        [44:0]   _zz_210;
  reg        [44:0]   _zz_211;
  reg        [44:0]   _zz_212;
  reg        [44:0]   _zz_213;
  reg        [44:0]   _zz_214;
  reg        [44:0]   _zz_215;
  reg        [47:0]   _zz_216;
  reg        [47:0]   _zz_217;
  reg        [47:0]   _zz_218;
  reg        [47:0]   _zz_219;
  reg        [47:0]   _zz_220;
  reg        [47:0]   _zz_221;
  reg        [47:0]   _zz_222;
  reg        [47:0]   _zz_223;
  reg        [47:0]   _zz_224;
  reg        [47:0]   _zz_225;
  reg        [47:0]   _zz_226;
  reg        [47:0]   _zz_227;
  reg        [47:0]   _zz_228;
  reg        [47:0]   _zz_229;
  reg        [47:0]   _zz_230;
  reg        [47:0]   _zz_231;
  reg        [47:0]   _zz_232;
  reg        [47:0]   _zz_233;
  reg        [47:0]   _zz_234;
  reg        [47:0]   _zz_235;
  reg        [47:0]   _zz_236;
  reg        [47:0]   _zz_237;
  reg        [47:0]   _zz_238;
  reg        [47:0]   _zz_239;
  reg        [47:0]   _zz_240;
  reg        [47:0]   _zz_241;
  reg        [47:0]   _zz_242;
  reg        [47:0]   _zz_243;
  reg        [47:0]   _zz_244;
  reg        [47:0]   _zz_245;
  reg        [47:0]   _zz_246;
  reg        [47:0]   _zz_247;
  reg        [47:0]   _zz_248;
  reg        [47:0]   _zz_249;
  reg        [47:0]   _zz_250;
  reg        [47:0]   _zz_251;
  reg        [47:0]   _zz_252;
  reg        [47:0]   _zz_253;
  reg        [47:0]   _zz_254;
  reg        [47:0]   _zz_255;
  reg        [47:0]   _zz_256;
  reg        [47:0]   _zz_257;
  reg        [47:0]   _zz_258;
  reg        [47:0]   _zz_259;
  reg        [47:0]   _zz_260;
  reg        [47:0]   _zz_261;
  reg        [47:0]   _zz_262;
  reg        [47:0]   _zz_263;
  reg        [47:0]   _zz_264;
  reg        [47:0]   _zz_265;
  reg        [47:0]   _zz_266;
  reg        [47:0]   _zz_267;
  reg        [47:0]   _zz_268;
  reg        [47:0]   _zz_269;
  reg        [47:0]   _zz_270;
  reg        [47:0]   _zz_271;
  reg        [47:0]   _zz_272;
  reg        [47:0]   _zz_273;
  reg        [47:0]   _zz_274;
  reg        [47:0]   _zz_275;
  reg        [47:0]   _zz_276;
  reg        [47:0]   _zz_277;
  reg        [47:0]   _zz_278;
  reg        [47:0]   _zz_279;
  reg        [47:0]   _zz_280;
  reg        [47:0]   _zz_281;
  reg        [47:0]   _zz_282;
  reg        [47:0]   _zz_283;
  reg        [47:0]   _zz_284;
  reg        [47:0]   _zz_285;
  reg        [47:0]   _zz_286;
  reg        [47:0]   _zz_287;
  reg        [47:0]   _zz_288;

  assign _zz_289 = {{3{_zz_145[44]}}, _zz_145};
  assign _zz_290 = {{3{_zz_146[44]}}, _zz_146};
  assign _zz_291 = {{3{_zz_147[44]}}, _zz_147};
  assign _zz_292 = {{3{_zz_148[44]}}, _zz_148};
  assign _zz_293 = {{3{_zz_149[44]}}, _zz_149};
  assign _zz_294 = {{3{_zz_150[44]}}, _zz_150};
  assign _zz_295 = {{3{_zz_151[44]}}, _zz_151};
  assign _zz_296 = {{3{_zz_152[44]}}, _zz_152};
  assign _zz_297 = {{3{_zz_153[44]}}, _zz_153};
  assign _zz_298 = {{3{_zz_154[44]}}, _zz_154};
  assign _zz_299 = {{3{_zz_155[44]}}, _zz_155};
  assign _zz_300 = {{3{_zz_156[44]}}, _zz_156};
  assign _zz_301 = {{3{_zz_157[44]}}, _zz_157};
  assign _zz_302 = {{3{_zz_158[44]}}, _zz_158};
  assign _zz_303 = {{3{_zz_159[44]}}, _zz_159};
  assign _zz_304 = {{3{_zz_160[44]}}, _zz_160};
  assign _zz_305 = {{3{_zz_161[44]}}, _zz_161};
  assign _zz_306 = {{3{_zz_162[44]}}, _zz_162};
  assign _zz_307 = {{3{_zz_163[44]}}, _zz_163};
  assign _zz_308 = {{3{_zz_164[44]}}, _zz_164};
  assign _zz_309 = {{3{_zz_165[44]}}, _zz_165};
  assign _zz_310 = {{3{_zz_166[44]}}, _zz_166};
  assign _zz_311 = {{3{_zz_167[44]}}, _zz_167};
  assign _zz_312 = {{3{_zz_168[44]}}, _zz_168};
  assign _zz_313 = {{3{_zz_169[44]}}, _zz_169};
  assign _zz_314 = {{3{_zz_170[44]}}, _zz_170};
  assign _zz_315 = {{3{_zz_171[44]}}, _zz_171};
  assign _zz_316 = {{3{_zz_172[44]}}, _zz_172};
  assign _zz_317 = {{3{_zz_173[44]}}, _zz_173};
  assign _zz_318 = {{3{_zz_174[44]}}, _zz_174};
  assign _zz_319 = {{3{_zz_175[44]}}, _zz_175};
  assign _zz_320 = {{3{_zz_176[44]}}, _zz_176};
  assign _zz_321 = {{3{_zz_177[44]}}, _zz_177};
  assign _zz_322 = {{3{_zz_178[44]}}, _zz_178};
  assign _zz_323 = {{3{_zz_179[44]}}, _zz_179};
  assign _zz_324 = {{3{_zz_180[44]}}, _zz_180};
  assign _zz_325 = {{3{_zz_181[44]}}, _zz_181};
  assign _zz_326 = {{3{_zz_182[44]}}, _zz_182};
  assign _zz_327 = {{3{_zz_183[44]}}, _zz_183};
  assign _zz_328 = {{3{_zz_184[44]}}, _zz_184};
  assign _zz_329 = {{3{_zz_185[44]}}, _zz_185};
  assign _zz_330 = {{3{_zz_186[44]}}, _zz_186};
  assign _zz_331 = {{3{_zz_187[44]}}, _zz_187};
  assign _zz_332 = {{3{_zz_188[44]}}, _zz_188};
  assign _zz_333 = {{3{_zz_189[44]}}, _zz_189};
  assign _zz_334 = {{3{_zz_190[44]}}, _zz_190};
  assign _zz_335 = {{3{_zz_191[44]}}, _zz_191};
  assign _zz_336 = {{3{_zz_192[44]}}, _zz_192};
  assign _zz_337 = {{3{_zz_193[44]}}, _zz_193};
  assign _zz_338 = {{3{_zz_194[44]}}, _zz_194};
  assign _zz_339 = {{3{_zz_195[44]}}, _zz_195};
  assign _zz_340 = {{3{_zz_196[44]}}, _zz_196};
  assign _zz_341 = {{3{_zz_197[44]}}, _zz_197};
  assign _zz_342 = {{3{_zz_198[44]}}, _zz_198};
  assign _zz_343 = {{3{_zz_199[44]}}, _zz_199};
  assign _zz_344 = {{3{_zz_200[44]}}, _zz_200};
  assign _zz_345 = {{3{_zz_201[44]}}, _zz_201};
  assign _zz_346 = {{3{_zz_202[44]}}, _zz_202};
  assign _zz_347 = {{3{_zz_203[44]}}, _zz_203};
  assign _zz_348 = {{3{_zz_204[44]}}, _zz_204};
  assign _zz_349 = {{3{_zz_205[44]}}, _zz_205};
  assign _zz_350 = {{3{_zz_206[44]}}, _zz_206};
  assign _zz_351 = {{3{_zz_207[44]}}, _zz_207};
  assign _zz_352 = {{3{_zz_208[44]}}, _zz_208};
  assign _zz_353 = {{3{_zz_209[44]}}, _zz_209};
  assign _zz_354 = {{3{_zz_210[44]}}, _zz_210};
  assign _zz_355 = {{3{_zz_211[44]}}, _zz_211};
  assign _zz_356 = {{3{_zz_212[44]}}, _zz_212};
  assign _zz_357 = {{3{_zz_213[44]}}, _zz_213};
  assign _zz_358 = {{3{_zz_214[44]}}, _zz_214};
  assign _zz_359 = {{3{_zz_215[44]}}, _zz_215};
  assign weightWires_0 = 18'h001a1;
  assign weightWires_1 = 18'h00218;
  assign weightWires_2 = 18'h00213;
  assign weightWires_3 = 18'h0019c;
  assign weightWires_4 = 18'h0023d;
  assign weightWires_5 = 18'h001f4;
  assign weightWires_6 = 18'h001dd;
  assign weightWires_7 = 18'h001d5;
  assign weightWires_8 = 18'h0020d;
  assign weightWires_9 = 18'h00253;
  assign weightWires_10 = 18'h00233;
  assign weightWires_11 = 18'h0019c;
  assign weightWires_12 = 18'h0019b;
  assign weightWires_13 = 18'h00215;
  assign weightWires_14 = 18'h00253;
  assign weightWires_15 = 18'h001a8;
  assign weightWires_16 = 18'h00239;
  assign weightWires_17 = 18'h001f0;
  assign weightWires_18 = 18'h001a6;
  assign weightWires_19 = 18'h001fb;
  assign weightWires_20 = 18'h001ed;
  assign weightWires_21 = 18'h001b2;
  assign weightWires_22 = 18'h00196;
  assign weightWires_23 = 18'h001dc;
  assign weightWires_24 = 18'h0021a;
  assign weightWires_25 = 18'h001be;
  assign weightWires_26 = 18'h00231;
  assign weightWires_27 = 18'h001e8;
  assign weightWires_28 = 18'h00227;
  assign weightWires_29 = 18'h001ed;
  assign weightWires_30 = 18'h0024d;
  assign weightWires_31 = 18'h00241;
  assign weightWires_32 = 18'h00195;
  assign weightWires_33 = 18'h001c9;
  assign weightWires_34 = 18'h0023d;
  assign weightWires_35 = 18'h00255;
  assign weightWires_36 = 18'h001e5;
  assign weightWires_37 = 18'h0024a;
  assign weightWires_38 = 18'h001bf;
  assign weightWires_39 = 18'h001e3;
  assign weightWires_40 = 18'h001d9;
  assign weightWires_41 = 18'h00211;
  assign weightWires_42 = 18'h001b7;
  assign weightWires_43 = 18'h00256;
  assign weightWires_44 = 18'h0022e;
  assign weightWires_45 = 18'h001da;
  assign weightWires_46 = 18'h00194;
  assign weightWires_47 = 18'h001cb;
  assign weightWires_48 = 18'h0023b;
  assign weightWires_49 = 18'h001ce;
  assign weightWires_50 = 18'h0023c;
  assign weightWires_51 = 18'h0024d;
  assign weightWires_52 = 18'h001ac;
  assign weightWires_53 = 18'h001f3;
  assign weightWires_54 = 18'h00239;
  assign weightWires_55 = 18'h0024e;
  assign weightWires_56 = 18'h00202;
  assign weightWires_57 = 18'h00235;
  assign weightWires_58 = 18'h0022a;
  assign weightWires_59 = 18'h001c4;
  assign weightWires_60 = 18'h00216;
  assign weightWires_61 = 18'h0020e;
  assign weightWires_62 = 18'h001c3;
  assign weightWires_63 = 18'h001b8;
  assign weightWires_64 = 18'h001d3;
  assign weightWires_65 = 18'h00242;
  assign weightWires_66 = 18'h0020d;
  assign weightWires_67 = 18'h001e6;
  assign weightWires_68 = 18'h00214;
  assign weightWires_69 = 18'h001a1;
  assign weightWires_70 = 18'h00198;
  assign weightWires_71 = 18'h001b2;
  assign inputZERO = 27'h0;
  assign io_dataOut = _zz_288;
  always @ (posedge clk) begin
    io_dataIn_regNext <= io_dataIn;
    _zz_1 <= io_dataIn_regNext;
    _zz_144 <= ($signed(weightWires_0) * $signed(_zz_1));
    _zz_216 <= {{3{_zz_144[44]}}, _zz_144};
    _zz_2 <= _zz_1;
    _zz_3 <= _zz_2;
    _zz_145 <= ($signed(weightWires_1) * $signed(_zz_3));
    _zz_217 <= ($signed(_zz_216) + $signed(_zz_289));
    _zz_4 <= _zz_3;
    _zz_5 <= _zz_4;
    _zz_146 <= ($signed(weightWires_2) * $signed(_zz_5));
    _zz_218 <= ($signed(_zz_217) + $signed(_zz_290));
    _zz_6 <= _zz_5;
    _zz_7 <= _zz_6;
    _zz_147 <= ($signed(weightWires_3) * $signed(_zz_7));
    _zz_219 <= ($signed(_zz_218) + $signed(_zz_291));
    _zz_8 <= _zz_7;
    _zz_9 <= _zz_8;
    _zz_148 <= ($signed(weightWires_4) * $signed(_zz_9));
    _zz_220 <= ($signed(_zz_219) + $signed(_zz_292));
    _zz_10 <= _zz_9;
    _zz_11 <= _zz_10;
    _zz_149 <= ($signed(weightWires_5) * $signed(_zz_11));
    _zz_221 <= ($signed(_zz_220) + $signed(_zz_293));
    _zz_12 <= _zz_11;
    _zz_13 <= _zz_12;
    _zz_150 <= ($signed(weightWires_6) * $signed(_zz_13));
    _zz_222 <= ($signed(_zz_221) + $signed(_zz_294));
    _zz_14 <= _zz_13;
    _zz_15 <= _zz_14;
    _zz_151 <= ($signed(weightWires_7) * $signed(_zz_15));
    _zz_223 <= ($signed(_zz_222) + $signed(_zz_295));
    _zz_16 <= _zz_15;
    _zz_17 <= _zz_16;
    _zz_152 <= ($signed(weightWires_8) * $signed(_zz_17));
    _zz_224 <= ($signed(_zz_223) + $signed(_zz_296));
    _zz_18 <= _zz_17;
    _zz_19 <= _zz_18;
    _zz_153 <= ($signed(weightWires_9) * $signed(_zz_19));
    _zz_225 <= ($signed(_zz_224) + $signed(_zz_297));
    _zz_20 <= _zz_19;
    _zz_21 <= _zz_20;
    _zz_154 <= ($signed(weightWires_10) * $signed(_zz_21));
    _zz_226 <= ($signed(_zz_225) + $signed(_zz_298));
    _zz_22 <= _zz_21;
    _zz_23 <= _zz_22;
    _zz_155 <= ($signed(weightWires_11) * $signed(_zz_23));
    _zz_227 <= ($signed(_zz_226) + $signed(_zz_299));
    _zz_24 <= _zz_23;
    _zz_25 <= _zz_24;
    _zz_156 <= ($signed(weightWires_12) * $signed(_zz_25));
    _zz_228 <= ($signed(_zz_227) + $signed(_zz_300));
    _zz_26 <= _zz_25;
    _zz_27 <= _zz_26;
    _zz_157 <= ($signed(weightWires_13) * $signed(_zz_27));
    _zz_229 <= ($signed(_zz_228) + $signed(_zz_301));
    _zz_28 <= _zz_27;
    _zz_29 <= _zz_28;
    _zz_158 <= ($signed(weightWires_14) * $signed(_zz_29));
    _zz_230 <= ($signed(_zz_229) + $signed(_zz_302));
    _zz_30 <= _zz_29;
    _zz_31 <= _zz_30;
    _zz_159 <= ($signed(weightWires_15) * $signed(_zz_31));
    _zz_231 <= ($signed(_zz_230) + $signed(_zz_303));
    _zz_32 <= _zz_31;
    _zz_33 <= _zz_32;
    _zz_160 <= ($signed(weightWires_16) * $signed(_zz_33));
    _zz_232 <= ($signed(_zz_231) + $signed(_zz_304));
    _zz_34 <= _zz_33;
    _zz_35 <= _zz_34;
    _zz_161 <= ($signed(weightWires_17) * $signed(_zz_35));
    _zz_233 <= ($signed(_zz_232) + $signed(_zz_305));
    _zz_36 <= _zz_35;
    _zz_37 <= _zz_36;
    _zz_162 <= ($signed(weightWires_18) * $signed(_zz_37));
    _zz_234 <= ($signed(_zz_233) + $signed(_zz_306));
    _zz_38 <= _zz_37;
    _zz_39 <= _zz_38;
    _zz_163 <= ($signed(weightWires_19) * $signed(_zz_39));
    _zz_235 <= ($signed(_zz_234) + $signed(_zz_307));
    _zz_40 <= _zz_39;
    _zz_41 <= _zz_40;
    _zz_164 <= ($signed(weightWires_20) * $signed(_zz_41));
    _zz_236 <= ($signed(_zz_235) + $signed(_zz_308));
    _zz_42 <= _zz_41;
    _zz_43 <= _zz_42;
    _zz_165 <= ($signed(weightWires_21) * $signed(_zz_43));
    _zz_237 <= ($signed(_zz_236) + $signed(_zz_309));
    _zz_44 <= _zz_43;
    _zz_45 <= _zz_44;
    _zz_166 <= ($signed(weightWires_22) * $signed(_zz_45));
    _zz_238 <= ($signed(_zz_237) + $signed(_zz_310));
    _zz_46 <= _zz_45;
    _zz_47 <= _zz_46;
    _zz_167 <= ($signed(weightWires_23) * $signed(_zz_47));
    _zz_239 <= ($signed(_zz_238) + $signed(_zz_311));
    _zz_48 <= _zz_47;
    _zz_49 <= _zz_48;
    _zz_168 <= ($signed(weightWires_24) * $signed(_zz_49));
    _zz_240 <= ($signed(_zz_239) + $signed(_zz_312));
    _zz_50 <= _zz_49;
    _zz_51 <= _zz_50;
    _zz_169 <= ($signed(weightWires_25) * $signed(_zz_51));
    _zz_241 <= ($signed(_zz_240) + $signed(_zz_313));
    _zz_52 <= _zz_51;
    _zz_53 <= _zz_52;
    _zz_170 <= ($signed(weightWires_26) * $signed(_zz_53));
    _zz_242 <= ($signed(_zz_241) + $signed(_zz_314));
    _zz_54 <= _zz_53;
    _zz_55 <= _zz_54;
    _zz_171 <= ($signed(weightWires_27) * $signed(_zz_55));
    _zz_243 <= ($signed(_zz_242) + $signed(_zz_315));
    _zz_56 <= _zz_55;
    _zz_57 <= _zz_56;
    _zz_172 <= ($signed(weightWires_28) * $signed(_zz_57));
    _zz_244 <= ($signed(_zz_243) + $signed(_zz_316));
    _zz_58 <= _zz_57;
    _zz_59 <= _zz_58;
    _zz_173 <= ($signed(weightWires_29) * $signed(_zz_59));
    _zz_245 <= ($signed(_zz_244) + $signed(_zz_317));
    _zz_60 <= _zz_59;
    _zz_61 <= _zz_60;
    _zz_174 <= ($signed(weightWires_30) * $signed(_zz_61));
    _zz_246 <= ($signed(_zz_245) + $signed(_zz_318));
    _zz_62 <= _zz_61;
    _zz_63 <= _zz_62;
    _zz_175 <= ($signed(weightWires_31) * $signed(_zz_63));
    _zz_247 <= ($signed(_zz_246) + $signed(_zz_319));
    _zz_64 <= _zz_63;
    _zz_65 <= _zz_64;
    _zz_176 <= ($signed(weightWires_32) * $signed(_zz_65));
    _zz_248 <= ($signed(_zz_247) + $signed(_zz_320));
    _zz_66 <= _zz_65;
    _zz_67 <= _zz_66;
    _zz_177 <= ($signed(weightWires_33) * $signed(_zz_67));
    _zz_249 <= ($signed(_zz_248) + $signed(_zz_321));
    _zz_68 <= _zz_67;
    _zz_69 <= _zz_68;
    _zz_178 <= ($signed(weightWires_34) * $signed(_zz_69));
    _zz_250 <= ($signed(_zz_249) + $signed(_zz_322));
    _zz_70 <= _zz_69;
    _zz_71 <= _zz_70;
    _zz_179 <= ($signed(weightWires_35) * $signed(_zz_71));
    _zz_251 <= ($signed(_zz_250) + $signed(_zz_323));
    _zz_72 <= _zz_71;
    _zz_73 <= _zz_72;
    _zz_180 <= ($signed(weightWires_36) * $signed(_zz_73));
    _zz_252 <= ($signed(_zz_251) + $signed(_zz_324));
    _zz_74 <= _zz_73;
    _zz_75 <= _zz_74;
    _zz_181 <= ($signed(weightWires_37) * $signed(_zz_75));
    _zz_253 <= ($signed(_zz_252) + $signed(_zz_325));
    _zz_76 <= _zz_75;
    _zz_77 <= _zz_76;
    _zz_182 <= ($signed(weightWires_38) * $signed(_zz_77));
    _zz_254 <= ($signed(_zz_253) + $signed(_zz_326));
    _zz_78 <= _zz_77;
    _zz_79 <= _zz_78;
    _zz_183 <= ($signed(weightWires_39) * $signed(_zz_79));
    _zz_255 <= ($signed(_zz_254) + $signed(_zz_327));
    _zz_80 <= _zz_79;
    _zz_81 <= _zz_80;
    _zz_184 <= ($signed(weightWires_40) * $signed(_zz_81));
    _zz_256 <= ($signed(_zz_255) + $signed(_zz_328));
    _zz_82 <= _zz_81;
    _zz_83 <= _zz_82;
    _zz_185 <= ($signed(weightWires_41) * $signed(_zz_83));
    _zz_257 <= ($signed(_zz_256) + $signed(_zz_329));
    _zz_84 <= _zz_83;
    _zz_85 <= _zz_84;
    _zz_186 <= ($signed(weightWires_42) * $signed(_zz_85));
    _zz_258 <= ($signed(_zz_257) + $signed(_zz_330));
    _zz_86 <= _zz_85;
    _zz_87 <= _zz_86;
    _zz_187 <= ($signed(weightWires_43) * $signed(_zz_87));
    _zz_259 <= ($signed(_zz_258) + $signed(_zz_331));
    _zz_88 <= _zz_87;
    _zz_89 <= _zz_88;
    _zz_188 <= ($signed(weightWires_44) * $signed(_zz_89));
    _zz_260 <= ($signed(_zz_259) + $signed(_zz_332));
    _zz_90 <= _zz_89;
    _zz_91 <= _zz_90;
    _zz_189 <= ($signed(weightWires_45) * $signed(_zz_91));
    _zz_261 <= ($signed(_zz_260) + $signed(_zz_333));
    _zz_92 <= _zz_91;
    _zz_93 <= _zz_92;
    _zz_190 <= ($signed(weightWires_46) * $signed(_zz_93));
    _zz_262 <= ($signed(_zz_261) + $signed(_zz_334));
    _zz_94 <= _zz_93;
    _zz_95 <= _zz_94;
    _zz_191 <= ($signed(weightWires_47) * $signed(_zz_95));
    _zz_263 <= ($signed(_zz_262) + $signed(_zz_335));
    _zz_96 <= _zz_95;
    _zz_97 <= _zz_96;
    _zz_192 <= ($signed(weightWires_48) * $signed(_zz_97));
    _zz_264 <= ($signed(_zz_263) + $signed(_zz_336));
    _zz_98 <= _zz_97;
    _zz_99 <= _zz_98;
    _zz_193 <= ($signed(weightWires_49) * $signed(_zz_99));
    _zz_265 <= ($signed(_zz_264) + $signed(_zz_337));
    _zz_100 <= _zz_99;
    _zz_101 <= _zz_100;
    _zz_194 <= ($signed(weightWires_50) * $signed(_zz_101));
    _zz_266 <= ($signed(_zz_265) + $signed(_zz_338));
    _zz_102 <= _zz_101;
    _zz_103 <= _zz_102;
    _zz_195 <= ($signed(weightWires_51) * $signed(_zz_103));
    _zz_267 <= ($signed(_zz_266) + $signed(_zz_339));
    _zz_104 <= _zz_103;
    _zz_105 <= _zz_104;
    _zz_196 <= ($signed(weightWires_52) * $signed(_zz_105));
    _zz_268 <= ($signed(_zz_267) + $signed(_zz_340));
    _zz_106 <= _zz_105;
    _zz_107 <= _zz_106;
    _zz_197 <= ($signed(weightWires_53) * $signed(_zz_107));
    _zz_269 <= ($signed(_zz_268) + $signed(_zz_341));
    _zz_108 <= _zz_107;
    _zz_109 <= _zz_108;
    _zz_198 <= ($signed(weightWires_54) * $signed(_zz_109));
    _zz_270 <= ($signed(_zz_269) + $signed(_zz_342));
    _zz_110 <= _zz_109;
    _zz_111 <= _zz_110;
    _zz_199 <= ($signed(weightWires_55) * $signed(_zz_111));
    _zz_271 <= ($signed(_zz_270) + $signed(_zz_343));
    _zz_112 <= _zz_111;
    _zz_113 <= _zz_112;
    _zz_200 <= ($signed(weightWires_56) * $signed(_zz_113));
    _zz_272 <= ($signed(_zz_271) + $signed(_zz_344));
    _zz_114 <= _zz_113;
    _zz_115 <= _zz_114;
    _zz_201 <= ($signed(weightWires_57) * $signed(_zz_115));
    _zz_273 <= ($signed(_zz_272) + $signed(_zz_345));
    _zz_116 <= _zz_115;
    _zz_117 <= _zz_116;
    _zz_202 <= ($signed(weightWires_58) * $signed(_zz_117));
    _zz_274 <= ($signed(_zz_273) + $signed(_zz_346));
    _zz_118 <= _zz_117;
    _zz_119 <= _zz_118;
    _zz_203 <= ($signed(weightWires_59) * $signed(_zz_119));
    _zz_275 <= ($signed(_zz_274) + $signed(_zz_347));
    _zz_120 <= _zz_119;
    _zz_121 <= _zz_120;
    _zz_204 <= ($signed(weightWires_60) * $signed(_zz_121));
    _zz_276 <= ($signed(_zz_275) + $signed(_zz_348));
    _zz_122 <= _zz_121;
    _zz_123 <= _zz_122;
    _zz_205 <= ($signed(weightWires_61) * $signed(_zz_123));
    _zz_277 <= ($signed(_zz_276) + $signed(_zz_349));
    _zz_124 <= _zz_123;
    _zz_125 <= _zz_124;
    _zz_206 <= ($signed(weightWires_62) * $signed(_zz_125));
    _zz_278 <= ($signed(_zz_277) + $signed(_zz_350));
    _zz_126 <= _zz_125;
    _zz_127 <= _zz_126;
    _zz_207 <= ($signed(weightWires_63) * $signed(_zz_127));
    _zz_279 <= ($signed(_zz_278) + $signed(_zz_351));
    _zz_128 <= _zz_127;
    _zz_129 <= _zz_128;
    _zz_208 <= ($signed(weightWires_64) * $signed(_zz_129));
    _zz_280 <= ($signed(_zz_279) + $signed(_zz_352));
    _zz_130 <= _zz_129;
    _zz_131 <= _zz_130;
    _zz_209 <= ($signed(weightWires_65) * $signed(_zz_131));
    _zz_281 <= ($signed(_zz_280) + $signed(_zz_353));
    _zz_132 <= _zz_131;
    _zz_133 <= _zz_132;
    _zz_210 <= ($signed(weightWires_66) * $signed(_zz_133));
    _zz_282 <= ($signed(_zz_281) + $signed(_zz_354));
    _zz_134 <= _zz_133;
    _zz_135 <= _zz_134;
    _zz_211 <= ($signed(weightWires_67) * $signed(_zz_135));
    _zz_283 <= ($signed(_zz_282) + $signed(_zz_355));
    _zz_136 <= _zz_135;
    _zz_137 <= _zz_136;
    _zz_212 <= ($signed(weightWires_68) * $signed(_zz_137));
    _zz_284 <= ($signed(_zz_283) + $signed(_zz_356));
    _zz_138 <= _zz_137;
    _zz_139 <= _zz_138;
    _zz_213 <= ($signed(weightWires_69) * $signed(_zz_139));
    _zz_285 <= ($signed(_zz_284) + $signed(_zz_357));
    _zz_140 <= _zz_139;
    _zz_141 <= _zz_140;
    _zz_214 <= ($signed(weightWires_70) * $signed(_zz_141));
    _zz_286 <= ($signed(_zz_285) + $signed(_zz_358));
    _zz_142 <= _zz_141;
    _zz_143 <= _zz_142;
    _zz_215 <= ($signed(weightWires_71) * $signed(_zz_143));
    _zz_287 <= ($signed(_zz_286) + $signed(_zz_359));
    _zz_288 <= _zz_287;
  end


endmodule
