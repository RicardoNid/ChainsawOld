// lsfan
// 2020��11��30��

module regs_ifid (
	input logic clk,
	input logic rstn,
	output logic out
);
  
  f
  
  endmodule 