// Generator : SpinalHDL v1.4.2    git head : 804c7bd7b7feaddcc1d25ecef6c208fd5f776f79
// Component : Calc
// Git hash  : 9bc1f6abee76360b92dc957c4d115e31fb5afd89



module Calc (
  input               io_inputDataIn_valid,
  output              io_inputDataIn_ready,
  input      [7:0]    io_inputDataIn_payload_0,
  input      [7:0]    io_inputDataIn_payload_1,
  input      [7:0]    io_inputDataIn_payload_2,
  input      [7:0]    io_inputDataIn_payload_3,
  input      [7:0]    io_inputDataIn_payload_4,
  input      [7:0]    io_inputDataIn_payload_5,
  input      [7:0]    io_inputDataIn_payload_6,
  input      [7:0]    io_inputDataIn_payload_7,
  input      [7:0]    io_inputDataIn_payload_8,
  input      [7:0]    io_inputDataIn_payload_9,
  input      [7:0]    io_inputDataIn_payload_10,
  input      [7:0]    io_inputDataIn_payload_11,
  input      [7:0]    io_inputDataIn_payload_12,
  input      [7:0]    io_inputDataIn_payload_13,
  input      [7:0]    io_inputDataIn_payload_14,
  input      [7:0]    io_inputDataIn_payload_15,
  input               io_weightDataIn_valid,
  output              io_weightDataIn_ready,
  input      [7:0]    io_weightDataIn_payload_0_0,
  input      [7:0]    io_weightDataIn_payload_0_1,
  input      [7:0]    io_weightDataIn_payload_0_2,
  input      [7:0]    io_weightDataIn_payload_0_3,
  input      [7:0]    io_weightDataIn_payload_0_4,
  input      [7:0]    io_weightDataIn_payload_0_5,
  input      [7:0]    io_weightDataIn_payload_0_6,
  input      [7:0]    io_weightDataIn_payload_0_7,
  input      [7:0]    io_weightDataIn_payload_0_8,
  input      [7:0]    io_weightDataIn_payload_0_9,
  input      [7:0]    io_weightDataIn_payload_0_10,
  input      [7:0]    io_weightDataIn_payload_0_11,
  input      [7:0]    io_weightDataIn_payload_0_12,
  input      [7:0]    io_weightDataIn_payload_0_13,
  input      [7:0]    io_weightDataIn_payload_0_14,
  input      [7:0]    io_weightDataIn_payload_0_15,
  input      [7:0]    io_weightDataIn_payload_1_0,
  input      [7:0]    io_weightDataIn_payload_1_1,
  input      [7:0]    io_weightDataIn_payload_1_2,
  input      [7:0]    io_weightDataIn_payload_1_3,
  input      [7:0]    io_weightDataIn_payload_1_4,
  input      [7:0]    io_weightDataIn_payload_1_5,
  input      [7:0]    io_weightDataIn_payload_1_6,
  input      [7:0]    io_weightDataIn_payload_1_7,
  input      [7:0]    io_weightDataIn_payload_1_8,
  input      [7:0]    io_weightDataIn_payload_1_9,
  input      [7:0]    io_weightDataIn_payload_1_10,
  input      [7:0]    io_weightDataIn_payload_1_11,
  input      [7:0]    io_weightDataIn_payload_1_12,
  input      [7:0]    io_weightDataIn_payload_1_13,
  input      [7:0]    io_weightDataIn_payload_1_14,
  input      [7:0]    io_weightDataIn_payload_1_15,
  input      [7:0]    io_weightDataIn_payload_2_0,
  input      [7:0]    io_weightDataIn_payload_2_1,
  input      [7:0]    io_weightDataIn_payload_2_2,
  input      [7:0]    io_weightDataIn_payload_2_3,
  input      [7:0]    io_weightDataIn_payload_2_4,
  input      [7:0]    io_weightDataIn_payload_2_5,
  input      [7:0]    io_weightDataIn_payload_2_6,
  input      [7:0]    io_weightDataIn_payload_2_7,
  input      [7:0]    io_weightDataIn_payload_2_8,
  input      [7:0]    io_weightDataIn_payload_2_9,
  input      [7:0]    io_weightDataIn_payload_2_10,
  input      [7:0]    io_weightDataIn_payload_2_11,
  input      [7:0]    io_weightDataIn_payload_2_12,
  input      [7:0]    io_weightDataIn_payload_2_13,
  input      [7:0]    io_weightDataIn_payload_2_14,
  input      [7:0]    io_weightDataIn_payload_2_15,
  input      [7:0]    io_weightDataIn_payload_3_0,
  input      [7:0]    io_weightDataIn_payload_3_1,
  input      [7:0]    io_weightDataIn_payload_3_2,
  input      [7:0]    io_weightDataIn_payload_3_3,
  input      [7:0]    io_weightDataIn_payload_3_4,
  input      [7:0]    io_weightDataIn_payload_3_5,
  input      [7:0]    io_weightDataIn_payload_3_6,
  input      [7:0]    io_weightDataIn_payload_3_7,
  input      [7:0]    io_weightDataIn_payload_3_8,
  input      [7:0]    io_weightDataIn_payload_3_9,
  input      [7:0]    io_weightDataIn_payload_3_10,
  input      [7:0]    io_weightDataIn_payload_3_11,
  input      [7:0]    io_weightDataIn_payload_3_12,
  input      [7:0]    io_weightDataIn_payload_3_13,
  input      [7:0]    io_weightDataIn_payload_3_14,
  input      [7:0]    io_weightDataIn_payload_3_15,
  input      [7:0]    io_weightDataIn_payload_4_0,
  input      [7:0]    io_weightDataIn_payload_4_1,
  input      [7:0]    io_weightDataIn_payload_4_2,
  input      [7:0]    io_weightDataIn_payload_4_3,
  input      [7:0]    io_weightDataIn_payload_4_4,
  input      [7:0]    io_weightDataIn_payload_4_5,
  input      [7:0]    io_weightDataIn_payload_4_6,
  input      [7:0]    io_weightDataIn_payload_4_7,
  input      [7:0]    io_weightDataIn_payload_4_8,
  input      [7:0]    io_weightDataIn_payload_4_9,
  input      [7:0]    io_weightDataIn_payload_4_10,
  input      [7:0]    io_weightDataIn_payload_4_11,
  input      [7:0]    io_weightDataIn_payload_4_12,
  input      [7:0]    io_weightDataIn_payload_4_13,
  input      [7:0]    io_weightDataIn_payload_4_14,
  input      [7:0]    io_weightDataIn_payload_4_15,
  input      [7:0]    io_weightDataIn_payload_5_0,
  input      [7:0]    io_weightDataIn_payload_5_1,
  input      [7:0]    io_weightDataIn_payload_5_2,
  input      [7:0]    io_weightDataIn_payload_5_3,
  input      [7:0]    io_weightDataIn_payload_5_4,
  input      [7:0]    io_weightDataIn_payload_5_5,
  input      [7:0]    io_weightDataIn_payload_5_6,
  input      [7:0]    io_weightDataIn_payload_5_7,
  input      [7:0]    io_weightDataIn_payload_5_8,
  input      [7:0]    io_weightDataIn_payload_5_9,
  input      [7:0]    io_weightDataIn_payload_5_10,
  input      [7:0]    io_weightDataIn_payload_5_11,
  input      [7:0]    io_weightDataIn_payload_5_12,
  input      [7:0]    io_weightDataIn_payload_5_13,
  input      [7:0]    io_weightDataIn_payload_5_14,
  input      [7:0]    io_weightDataIn_payload_5_15,
  input      [7:0]    io_weightDataIn_payload_6_0,
  input      [7:0]    io_weightDataIn_payload_6_1,
  input      [7:0]    io_weightDataIn_payload_6_2,
  input      [7:0]    io_weightDataIn_payload_6_3,
  input      [7:0]    io_weightDataIn_payload_6_4,
  input      [7:0]    io_weightDataIn_payload_6_5,
  input      [7:0]    io_weightDataIn_payload_6_6,
  input      [7:0]    io_weightDataIn_payload_6_7,
  input      [7:0]    io_weightDataIn_payload_6_8,
  input      [7:0]    io_weightDataIn_payload_6_9,
  input      [7:0]    io_weightDataIn_payload_6_10,
  input      [7:0]    io_weightDataIn_payload_6_11,
  input      [7:0]    io_weightDataIn_payload_6_12,
  input      [7:0]    io_weightDataIn_payload_6_13,
  input      [7:0]    io_weightDataIn_payload_6_14,
  input      [7:0]    io_weightDataIn_payload_6_15,
  input      [7:0]    io_weightDataIn_payload_7_0,
  input      [7:0]    io_weightDataIn_payload_7_1,
  input      [7:0]    io_weightDataIn_payload_7_2,
  input      [7:0]    io_weightDataIn_payload_7_3,
  input      [7:0]    io_weightDataIn_payload_7_4,
  input      [7:0]    io_weightDataIn_payload_7_5,
  input      [7:0]    io_weightDataIn_payload_7_6,
  input      [7:0]    io_weightDataIn_payload_7_7,
  input      [7:0]    io_weightDataIn_payload_7_8,
  input      [7:0]    io_weightDataIn_payload_7_9,
  input      [7:0]    io_weightDataIn_payload_7_10,
  input      [7:0]    io_weightDataIn_payload_7_11,
  input      [7:0]    io_weightDataIn_payload_7_12,
  input      [7:0]    io_weightDataIn_payload_7_13,
  input      [7:0]    io_weightDataIn_payload_7_14,
  input      [7:0]    io_weightDataIn_payload_7_15,
  input      [7:0]    io_weightDataIn_payload_8_0,
  input      [7:0]    io_weightDataIn_payload_8_1,
  input      [7:0]    io_weightDataIn_payload_8_2,
  input      [7:0]    io_weightDataIn_payload_8_3,
  input      [7:0]    io_weightDataIn_payload_8_4,
  input      [7:0]    io_weightDataIn_payload_8_5,
  input      [7:0]    io_weightDataIn_payload_8_6,
  input      [7:0]    io_weightDataIn_payload_8_7,
  input      [7:0]    io_weightDataIn_payload_8_8,
  input      [7:0]    io_weightDataIn_payload_8_9,
  input      [7:0]    io_weightDataIn_payload_8_10,
  input      [7:0]    io_weightDataIn_payload_8_11,
  input      [7:0]    io_weightDataIn_payload_8_12,
  input      [7:0]    io_weightDataIn_payload_8_13,
  input      [7:0]    io_weightDataIn_payload_8_14,
  input      [7:0]    io_weightDataIn_payload_8_15,
  input      [7:0]    io_weightDataIn_payload_9_0,
  input      [7:0]    io_weightDataIn_payload_9_1,
  input      [7:0]    io_weightDataIn_payload_9_2,
  input      [7:0]    io_weightDataIn_payload_9_3,
  input      [7:0]    io_weightDataIn_payload_9_4,
  input      [7:0]    io_weightDataIn_payload_9_5,
  input      [7:0]    io_weightDataIn_payload_9_6,
  input      [7:0]    io_weightDataIn_payload_9_7,
  input      [7:0]    io_weightDataIn_payload_9_8,
  input      [7:0]    io_weightDataIn_payload_9_9,
  input      [7:0]    io_weightDataIn_payload_9_10,
  input      [7:0]    io_weightDataIn_payload_9_11,
  input      [7:0]    io_weightDataIn_payload_9_12,
  input      [7:0]    io_weightDataIn_payload_9_13,
  input      [7:0]    io_weightDataIn_payload_9_14,
  input      [7:0]    io_weightDataIn_payload_9_15,
  input      [7:0]    io_weightDataIn_payload_10_0,
  input      [7:0]    io_weightDataIn_payload_10_1,
  input      [7:0]    io_weightDataIn_payload_10_2,
  input      [7:0]    io_weightDataIn_payload_10_3,
  input      [7:0]    io_weightDataIn_payload_10_4,
  input      [7:0]    io_weightDataIn_payload_10_5,
  input      [7:0]    io_weightDataIn_payload_10_6,
  input      [7:0]    io_weightDataIn_payload_10_7,
  input      [7:0]    io_weightDataIn_payload_10_8,
  input      [7:0]    io_weightDataIn_payload_10_9,
  input      [7:0]    io_weightDataIn_payload_10_10,
  input      [7:0]    io_weightDataIn_payload_10_11,
  input      [7:0]    io_weightDataIn_payload_10_12,
  input      [7:0]    io_weightDataIn_payload_10_13,
  input      [7:0]    io_weightDataIn_payload_10_14,
  input      [7:0]    io_weightDataIn_payload_10_15,
  input      [7:0]    io_weightDataIn_payload_11_0,
  input      [7:0]    io_weightDataIn_payload_11_1,
  input      [7:0]    io_weightDataIn_payload_11_2,
  input      [7:0]    io_weightDataIn_payload_11_3,
  input      [7:0]    io_weightDataIn_payload_11_4,
  input      [7:0]    io_weightDataIn_payload_11_5,
  input      [7:0]    io_weightDataIn_payload_11_6,
  input      [7:0]    io_weightDataIn_payload_11_7,
  input      [7:0]    io_weightDataIn_payload_11_8,
  input      [7:0]    io_weightDataIn_payload_11_9,
  input      [7:0]    io_weightDataIn_payload_11_10,
  input      [7:0]    io_weightDataIn_payload_11_11,
  input      [7:0]    io_weightDataIn_payload_11_12,
  input      [7:0]    io_weightDataIn_payload_11_13,
  input      [7:0]    io_weightDataIn_payload_11_14,
  input      [7:0]    io_weightDataIn_payload_11_15,
  input      [7:0]    io_weightDataIn_payload_12_0,
  input      [7:0]    io_weightDataIn_payload_12_1,
  input      [7:0]    io_weightDataIn_payload_12_2,
  input      [7:0]    io_weightDataIn_payload_12_3,
  input      [7:0]    io_weightDataIn_payload_12_4,
  input      [7:0]    io_weightDataIn_payload_12_5,
  input      [7:0]    io_weightDataIn_payload_12_6,
  input      [7:0]    io_weightDataIn_payload_12_7,
  input      [7:0]    io_weightDataIn_payload_12_8,
  input      [7:0]    io_weightDataIn_payload_12_9,
  input      [7:0]    io_weightDataIn_payload_12_10,
  input      [7:0]    io_weightDataIn_payload_12_11,
  input      [7:0]    io_weightDataIn_payload_12_12,
  input      [7:0]    io_weightDataIn_payload_12_13,
  input      [7:0]    io_weightDataIn_payload_12_14,
  input      [7:0]    io_weightDataIn_payload_12_15,
  input      [7:0]    io_weightDataIn_payload_13_0,
  input      [7:0]    io_weightDataIn_payload_13_1,
  input      [7:0]    io_weightDataIn_payload_13_2,
  input      [7:0]    io_weightDataIn_payload_13_3,
  input      [7:0]    io_weightDataIn_payload_13_4,
  input      [7:0]    io_weightDataIn_payload_13_5,
  input      [7:0]    io_weightDataIn_payload_13_6,
  input      [7:0]    io_weightDataIn_payload_13_7,
  input      [7:0]    io_weightDataIn_payload_13_8,
  input      [7:0]    io_weightDataIn_payload_13_9,
  input      [7:0]    io_weightDataIn_payload_13_10,
  input      [7:0]    io_weightDataIn_payload_13_11,
  input      [7:0]    io_weightDataIn_payload_13_12,
  input      [7:0]    io_weightDataIn_payload_13_13,
  input      [7:0]    io_weightDataIn_payload_13_14,
  input      [7:0]    io_weightDataIn_payload_13_15,
  input      [7:0]    io_weightDataIn_payload_14_0,
  input      [7:0]    io_weightDataIn_payload_14_1,
  input      [7:0]    io_weightDataIn_payload_14_2,
  input      [7:0]    io_weightDataIn_payload_14_3,
  input      [7:0]    io_weightDataIn_payload_14_4,
  input      [7:0]    io_weightDataIn_payload_14_5,
  input      [7:0]    io_weightDataIn_payload_14_6,
  input      [7:0]    io_weightDataIn_payload_14_7,
  input      [7:0]    io_weightDataIn_payload_14_8,
  input      [7:0]    io_weightDataIn_payload_14_9,
  input      [7:0]    io_weightDataIn_payload_14_10,
  input      [7:0]    io_weightDataIn_payload_14_11,
  input      [7:0]    io_weightDataIn_payload_14_12,
  input      [7:0]    io_weightDataIn_payload_14_13,
  input      [7:0]    io_weightDataIn_payload_14_14,
  input      [7:0]    io_weightDataIn_payload_14_15,
  input      [7:0]    io_weightDataIn_payload_15_0,
  input      [7:0]    io_weightDataIn_payload_15_1,
  input      [7:0]    io_weightDataIn_payload_15_2,
  input      [7:0]    io_weightDataIn_payload_15_3,
  input      [7:0]    io_weightDataIn_payload_15_4,
  input      [7:0]    io_weightDataIn_payload_15_5,
  input      [7:0]    io_weightDataIn_payload_15_6,
  input      [7:0]    io_weightDataIn_payload_15_7,
  input      [7:0]    io_weightDataIn_payload_15_8,
  input      [7:0]    io_weightDataIn_payload_15_9,
  input      [7:0]    io_weightDataIn_payload_15_10,
  input      [7:0]    io_weightDataIn_payload_15_11,
  input      [7:0]    io_weightDataIn_payload_15_12,
  input      [7:0]    io_weightDataIn_payload_15_13,
  input      [7:0]    io_weightDataIn_payload_15_14,
  input      [7:0]    io_weightDataIn_payload_15_15,
  output              io_calc2write_1_valid,
  input               io_calc2write_1_ready,
  output     [7:0]    io_calc2write_1_payload_0,
  output     [7:0]    io_calc2write_1_payload_1,
  output     [7:0]    io_calc2write_1_payload_2,
  output     [7:0]    io_calc2write_1_payload_3,
  output     [7:0]    io_calc2write_1_payload_4,
  output     [7:0]    io_calc2write_1_payload_5,
  output     [7:0]    io_calc2write_1_payload_6,
  output     [7:0]    io_calc2write_1_payload_7,
  output     [7:0]    io_calc2write_1_payload_8,
  output     [7:0]    io_calc2write_1_payload_9,
  output     [7:0]    io_calc2write_1_payload_10,
  output     [7:0]    io_calc2write_1_payload_11,
  output     [7:0]    io_calc2write_1_payload_12,
  output     [7:0]    io_calc2write_1_payload_13,
  output     [7:0]    io_calc2write_1_payload_14,
  output     [7:0]    io_calc2write_1_payload_15,
  output     [19:0]   adderTrees_0_result,
  output     [19:0]   adderTrees_1_result,
  output     [19:0]   adderTrees_2_result,
  output     [19:0]   adderTrees_3_result,
  output     [19:0]   adderTrees_4_result,
  output     [19:0]   adderTrees_5_result,
  output     [19:0]   adderTrees_6_result,
  output     [19:0]   adderTrees_7_result,
  output     [19:0]   adderTrees_8_result,
  output     [19:0]   adderTrees_9_result,
  output     [19:0]   adderTrees_10_result,
  output     [19:0]   adderTrees_11_result,
  output     [19:0]   adderTrees_12_result,
  output     [19:0]   adderTrees_13_result,
  output     [19:0]   adderTrees_14_result,
  output     [19:0]   adderTrees_15_result,
  input               clk,
  input               reset
);
  wire       [0:0]    _zz_241;
  wire       [1:0]    _zz_242;
  wire       [21:0]   _zz_243;
  wire       [21:0]   _zz_244;
  wire       [21:0]   _zz_245;
  wire       [21:0]   _zz_246;
  wire       [21:0]   _zz_247;
  wire       [21:0]   _zz_248;
  wire       [21:0]   _zz_249;
  wire       [21:0]   _zz_250;
  wire       [21:0]   _zz_251;
  wire       [21:0]   _zz_252;
  wire       [21:0]   _zz_253;
  wire       [21:0]   _zz_254;
  wire       [21:0]   _zz_255;
  wire       [21:0]   _zz_256;
  wire       [21:0]   _zz_257;
  wire       [21:0]   _zz_258;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_0_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_1_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_2_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_3_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_4_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_5_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_6_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_7_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_8_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_9_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_10_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_11_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_12_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_13_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_14_15;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_0;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_1;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_2;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_3;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_4;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_5;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_6;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_7;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_8;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_9;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_10;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_11;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_12;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_13;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_14;
  (* use_dsp = "yes" *) wire       [15:0]   multRegs_15_15;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_1;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_2;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_3;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_4;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_5;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_6;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_7;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_8;
  reg        [16:0]   _zz_1_regNext;
  reg        [16:0]   _zz_2_regNext;
  reg        [16:0]   _zz_3_regNext;
  reg        [16:0]   _zz_4_regNext;
  reg        [16:0]   _zz_5_regNext;
  reg        [16:0]   _zz_6_regNext;
  reg        [16:0]   _zz_7_regNext;
  reg        [16:0]   _zz_8_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_9;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_10;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_11;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_12;
  reg        [17:0]   _zz_9_regNext;
  reg        [17:0]   _zz_10_regNext;
  reg        [17:0]   _zz_11_regNext;
  reg        [17:0]   _zz_12_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_13;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_14;
  reg        [18:0]   _zz_13_regNext;
  reg        [18:0]   _zz_14_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_15;
  reg        [19:0]   _zz_15_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_16;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_17;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_18;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_19;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_20;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_21;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_22;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_23;
  reg        [16:0]   _zz_16_regNext;
  reg        [16:0]   _zz_17_regNext;
  reg        [16:0]   _zz_18_regNext;
  reg        [16:0]   _zz_19_regNext;
  reg        [16:0]   _zz_20_regNext;
  reg        [16:0]   _zz_21_regNext;
  reg        [16:0]   _zz_22_regNext;
  reg        [16:0]   _zz_23_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_24;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_25;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_26;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_27;
  reg        [17:0]   _zz_24_regNext;
  reg        [17:0]   _zz_25_regNext;
  reg        [17:0]   _zz_26_regNext;
  reg        [17:0]   _zz_27_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_28;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_29;
  reg        [18:0]   _zz_28_regNext;
  reg        [18:0]   _zz_29_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_30;
  reg        [19:0]   _zz_30_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_31;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_32;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_33;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_34;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_35;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_36;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_37;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_38;
  reg        [16:0]   _zz_31_regNext;
  reg        [16:0]   _zz_32_regNext;
  reg        [16:0]   _zz_33_regNext;
  reg        [16:0]   _zz_34_regNext;
  reg        [16:0]   _zz_35_regNext;
  reg        [16:0]   _zz_36_regNext;
  reg        [16:0]   _zz_37_regNext;
  reg        [16:0]   _zz_38_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_39;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_40;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_41;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_42;
  reg        [17:0]   _zz_39_regNext;
  reg        [17:0]   _zz_40_regNext;
  reg        [17:0]   _zz_41_regNext;
  reg        [17:0]   _zz_42_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_43;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_44;
  reg        [18:0]   _zz_43_regNext;
  reg        [18:0]   _zz_44_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_45;
  reg        [19:0]   _zz_45_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_46;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_47;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_48;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_49;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_50;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_51;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_52;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_53;
  reg        [16:0]   _zz_46_regNext;
  reg        [16:0]   _zz_47_regNext;
  reg        [16:0]   _zz_48_regNext;
  reg        [16:0]   _zz_49_regNext;
  reg        [16:0]   _zz_50_regNext;
  reg        [16:0]   _zz_51_regNext;
  reg        [16:0]   _zz_52_regNext;
  reg        [16:0]   _zz_53_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_54;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_55;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_56;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_57;
  reg        [17:0]   _zz_54_regNext;
  reg        [17:0]   _zz_55_regNext;
  reg        [17:0]   _zz_56_regNext;
  reg        [17:0]   _zz_57_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_58;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_59;
  reg        [18:0]   _zz_58_regNext;
  reg        [18:0]   _zz_59_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_60;
  reg        [19:0]   _zz_60_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_61;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_62;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_63;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_64;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_65;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_66;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_67;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_68;
  reg        [16:0]   _zz_61_regNext;
  reg        [16:0]   _zz_62_regNext;
  reg        [16:0]   _zz_63_regNext;
  reg        [16:0]   _zz_64_regNext;
  reg        [16:0]   _zz_65_regNext;
  reg        [16:0]   _zz_66_regNext;
  reg        [16:0]   _zz_67_regNext;
  reg        [16:0]   _zz_68_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_69;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_70;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_71;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_72;
  reg        [17:0]   _zz_69_regNext;
  reg        [17:0]   _zz_70_regNext;
  reg        [17:0]   _zz_71_regNext;
  reg        [17:0]   _zz_72_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_73;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_74;
  reg        [18:0]   _zz_73_regNext;
  reg        [18:0]   _zz_74_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_75;
  reg        [19:0]   _zz_75_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_76;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_77;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_78;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_79;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_80;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_81;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_82;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_83;
  reg        [16:0]   _zz_76_regNext;
  reg        [16:0]   _zz_77_regNext;
  reg        [16:0]   _zz_78_regNext;
  reg        [16:0]   _zz_79_regNext;
  reg        [16:0]   _zz_80_regNext;
  reg        [16:0]   _zz_81_regNext;
  reg        [16:0]   _zz_82_regNext;
  reg        [16:0]   _zz_83_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_84;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_85;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_86;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_87;
  reg        [17:0]   _zz_84_regNext;
  reg        [17:0]   _zz_85_regNext;
  reg        [17:0]   _zz_86_regNext;
  reg        [17:0]   _zz_87_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_88;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_89;
  reg        [18:0]   _zz_88_regNext;
  reg        [18:0]   _zz_89_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_90;
  reg        [19:0]   _zz_90_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_91;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_92;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_93;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_94;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_95;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_96;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_97;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_98;
  reg        [16:0]   _zz_91_regNext;
  reg        [16:0]   _zz_92_regNext;
  reg        [16:0]   _zz_93_regNext;
  reg        [16:0]   _zz_94_regNext;
  reg        [16:0]   _zz_95_regNext;
  reg        [16:0]   _zz_96_regNext;
  reg        [16:0]   _zz_97_regNext;
  reg        [16:0]   _zz_98_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_99;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_100;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_101;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_102;
  reg        [17:0]   _zz_99_regNext;
  reg        [17:0]   _zz_100_regNext;
  reg        [17:0]   _zz_101_regNext;
  reg        [17:0]   _zz_102_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_103;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_104;
  reg        [18:0]   _zz_103_regNext;
  reg        [18:0]   _zz_104_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_105;
  reg        [19:0]   _zz_105_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_106;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_107;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_108;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_109;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_110;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_111;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_112;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_113;
  reg        [16:0]   _zz_106_regNext;
  reg        [16:0]   _zz_107_regNext;
  reg        [16:0]   _zz_108_regNext;
  reg        [16:0]   _zz_109_regNext;
  reg        [16:0]   _zz_110_regNext;
  reg        [16:0]   _zz_111_regNext;
  reg        [16:0]   _zz_112_regNext;
  reg        [16:0]   _zz_113_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_114;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_115;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_116;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_117;
  reg        [17:0]   _zz_114_regNext;
  reg        [17:0]   _zz_115_regNext;
  reg        [17:0]   _zz_116_regNext;
  reg        [17:0]   _zz_117_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_118;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_119;
  reg        [18:0]   _zz_118_regNext;
  reg        [18:0]   _zz_119_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_120;
  reg        [19:0]   _zz_120_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_121;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_122;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_123;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_124;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_125;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_126;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_127;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_128;
  reg        [16:0]   _zz_121_regNext;
  reg        [16:0]   _zz_122_regNext;
  reg        [16:0]   _zz_123_regNext;
  reg        [16:0]   _zz_124_regNext;
  reg        [16:0]   _zz_125_regNext;
  reg        [16:0]   _zz_126_regNext;
  reg        [16:0]   _zz_127_regNext;
  reg        [16:0]   _zz_128_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_129;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_130;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_131;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_132;
  reg        [17:0]   _zz_129_regNext;
  reg        [17:0]   _zz_130_regNext;
  reg        [17:0]   _zz_131_regNext;
  reg        [17:0]   _zz_132_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_133;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_134;
  reg        [18:0]   _zz_133_regNext;
  reg        [18:0]   _zz_134_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_135;
  reg        [19:0]   _zz_135_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_136;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_137;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_138;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_139;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_140;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_141;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_142;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_143;
  reg        [16:0]   _zz_136_regNext;
  reg        [16:0]   _zz_137_regNext;
  reg        [16:0]   _zz_138_regNext;
  reg        [16:0]   _zz_139_regNext;
  reg        [16:0]   _zz_140_regNext;
  reg        [16:0]   _zz_141_regNext;
  reg        [16:0]   _zz_142_regNext;
  reg        [16:0]   _zz_143_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_144;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_145;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_146;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_147;
  reg        [17:0]   _zz_144_regNext;
  reg        [17:0]   _zz_145_regNext;
  reg        [17:0]   _zz_146_regNext;
  reg        [17:0]   _zz_147_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_148;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_149;
  reg        [18:0]   _zz_148_regNext;
  reg        [18:0]   _zz_149_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_150;
  reg        [19:0]   _zz_150_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_151;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_152;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_153;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_154;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_155;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_156;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_157;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_158;
  reg        [16:0]   _zz_151_regNext;
  reg        [16:0]   _zz_152_regNext;
  reg        [16:0]   _zz_153_regNext;
  reg        [16:0]   _zz_154_regNext;
  reg        [16:0]   _zz_155_regNext;
  reg        [16:0]   _zz_156_regNext;
  reg        [16:0]   _zz_157_regNext;
  reg        [16:0]   _zz_158_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_159;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_160;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_161;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_162;
  reg        [17:0]   _zz_159_regNext;
  reg        [17:0]   _zz_160_regNext;
  reg        [17:0]   _zz_161_regNext;
  reg        [17:0]   _zz_162_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_163;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_164;
  reg        [18:0]   _zz_163_regNext;
  reg        [18:0]   _zz_164_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_165;
  reg        [19:0]   _zz_165_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_166;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_167;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_168;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_169;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_170;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_171;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_172;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_173;
  reg        [16:0]   _zz_166_regNext;
  reg        [16:0]   _zz_167_regNext;
  reg        [16:0]   _zz_168_regNext;
  reg        [16:0]   _zz_169_regNext;
  reg        [16:0]   _zz_170_regNext;
  reg        [16:0]   _zz_171_regNext;
  reg        [16:0]   _zz_172_regNext;
  reg        [16:0]   _zz_173_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_174;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_175;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_176;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_177;
  reg        [17:0]   _zz_174_regNext;
  reg        [17:0]   _zz_175_regNext;
  reg        [17:0]   _zz_176_regNext;
  reg        [17:0]   _zz_177_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_178;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_179;
  reg        [18:0]   _zz_178_regNext;
  reg        [18:0]   _zz_179_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_180;
  reg        [19:0]   _zz_180_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_181;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_182;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_183;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_184;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_185;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_186;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_187;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_188;
  reg        [16:0]   _zz_181_regNext;
  reg        [16:0]   _zz_182_regNext;
  reg        [16:0]   _zz_183_regNext;
  reg        [16:0]   _zz_184_regNext;
  reg        [16:0]   _zz_185_regNext;
  reg        [16:0]   _zz_186_regNext;
  reg        [16:0]   _zz_187_regNext;
  reg        [16:0]   _zz_188_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_189;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_190;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_191;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_192;
  reg        [17:0]   _zz_189_regNext;
  reg        [17:0]   _zz_190_regNext;
  reg        [17:0]   _zz_191_regNext;
  reg        [17:0]   _zz_192_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_193;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_194;
  reg        [18:0]   _zz_193_regNext;
  reg        [18:0]   _zz_194_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_195;
  reg        [19:0]   _zz_195_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_196;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_197;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_198;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_199;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_200;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_201;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_202;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_203;
  reg        [16:0]   _zz_196_regNext;
  reg        [16:0]   _zz_197_regNext;
  reg        [16:0]   _zz_198_regNext;
  reg        [16:0]   _zz_199_regNext;
  reg        [16:0]   _zz_200_regNext;
  reg        [16:0]   _zz_201_regNext;
  reg        [16:0]   _zz_202_regNext;
  reg        [16:0]   _zz_203_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_204;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_205;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_206;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_207;
  reg        [17:0]   _zz_204_regNext;
  reg        [17:0]   _zz_205_regNext;
  reg        [17:0]   _zz_206_regNext;
  reg        [17:0]   _zz_207_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_208;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_209;
  reg        [18:0]   _zz_208_regNext;
  reg        [18:0]   _zz_209_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_210;
  reg        [19:0]   _zz_210_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_211;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_212;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_213;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_214;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_215;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_216;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_217;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_218;
  reg        [16:0]   _zz_211_regNext;
  reg        [16:0]   _zz_212_regNext;
  reg        [16:0]   _zz_213_regNext;
  reg        [16:0]   _zz_214_regNext;
  reg        [16:0]   _zz_215_regNext;
  reg        [16:0]   _zz_216_regNext;
  reg        [16:0]   _zz_217_regNext;
  reg        [16:0]   _zz_218_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_219;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_220;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_221;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_222;
  reg        [17:0]   _zz_219_regNext;
  reg        [17:0]   _zz_220_regNext;
  reg        [17:0]   _zz_221_regNext;
  reg        [17:0]   _zz_222_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_223;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_224;
  reg        [18:0]   _zz_223_regNext;
  reg        [18:0]   _zz_224_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_225;
  reg        [19:0]   _zz_225_regNext;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_226;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_227;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_228;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_229;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_230;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_231;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_232;
  (* dont_touch = "yes" *) wire       [16:0]   _zz_233;
  reg        [16:0]   _zz_226_regNext;
  reg        [16:0]   _zz_227_regNext;
  reg        [16:0]   _zz_228_regNext;
  reg        [16:0]   _zz_229_regNext;
  reg        [16:0]   _zz_230_regNext;
  reg        [16:0]   _zz_231_regNext;
  reg        [16:0]   _zz_232_regNext;
  reg        [16:0]   _zz_233_regNext;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_234;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_235;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_236;
  (* dont_touch = "yes" *) wire       [17:0]   _zz_237;
  reg        [17:0]   _zz_234_regNext;
  reg        [17:0]   _zz_235_regNext;
  reg        [17:0]   _zz_236_regNext;
  reg        [17:0]   _zz_237_regNext;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_238;
  (* dont_touch = "yes" *) wire       [18:0]   _zz_239;
  reg        [18:0]   _zz_238_regNext;
  reg        [18:0]   _zz_239_regNext;
  (* dont_touch = "yes" *) wire       [19:0]   _zz_240;
  reg        [19:0]   _zz_240_regNext;
  reg        [21:0]   accRegs_0;
  reg        [21:0]   accRegs_1;
  reg        [21:0]   accRegs_2;
  reg        [21:0]   accRegs_3;
  reg        [21:0]   accRegs_4;
  reg        [21:0]   accRegs_5;
  reg        [21:0]   accRegs_6;
  reg        [21:0]   accRegs_7;
  reg        [21:0]   accRegs_8;
  reg        [21:0]   accRegs_9;
  reg        [21:0]   accRegs_10;
  reg        [21:0]   accRegs_11;
  reg        [21:0]   accRegs_12;
  reg        [21:0]   accRegs_13;
  reg        [21:0]   accRegs_14;
  reg        [21:0]   accRegs_15;
  reg                 validCounter_willIncrement;
  wire                validCounter_willClear;
  reg        [1:0]    validCounter_valueNext;
  reg        [1:0]    validCounter_value;
  wire                validCounter_willOverflowIfInc;
  wire                validCounter_willOverflow;
  reg                 validCounter_willOverflow_delay_1;
  reg                 validCounter_willOverflow_delay_2;
  reg                 validCounter_willOverflow_delay_3;
  reg                 validCounter_willOverflow_delay_4;
  reg                 validCounter_willOverflow_delay_5;

  assign _zz_241 = validCounter_willIncrement;
  assign _zz_242 = {1'd0, _zz_241};
  assign _zz_243 = {2'd0, adderTrees_0_result};
  assign _zz_244 = {2'd0, adderTrees_1_result};
  assign _zz_245 = {2'd0, adderTrees_2_result};
  assign _zz_246 = {2'd0, adderTrees_3_result};
  assign _zz_247 = {2'd0, adderTrees_4_result};
  assign _zz_248 = {2'd0, adderTrees_5_result};
  assign _zz_249 = {2'd0, adderTrees_6_result};
  assign _zz_250 = {2'd0, adderTrees_7_result};
  assign _zz_251 = {2'd0, adderTrees_8_result};
  assign _zz_252 = {2'd0, adderTrees_9_result};
  assign _zz_253 = {2'd0, adderTrees_10_result};
  assign _zz_254 = {2'd0, adderTrees_11_result};
  assign _zz_255 = {2'd0, adderTrees_12_result};
  assign _zz_256 = {2'd0, adderTrees_13_result};
  assign _zz_257 = {2'd0, adderTrees_14_result};
  assign _zz_258 = {2'd0, adderTrees_15_result};
  assign multRegs_0_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_0_0);
  assign multRegs_0_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_0_1);
  assign multRegs_0_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_0_2);
  assign multRegs_0_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_0_3);
  assign multRegs_0_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_0_4);
  assign multRegs_0_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_0_5);
  assign multRegs_0_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_0_6);
  assign multRegs_0_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_0_7);
  assign multRegs_0_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_0_8);
  assign multRegs_0_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_0_9);
  assign multRegs_0_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_0_10);
  assign multRegs_0_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_0_11);
  assign multRegs_0_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_0_12);
  assign multRegs_0_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_0_13);
  assign multRegs_0_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_0_14);
  assign multRegs_0_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_0_15);
  assign multRegs_1_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_1_0);
  assign multRegs_1_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_1_1);
  assign multRegs_1_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_1_2);
  assign multRegs_1_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_1_3);
  assign multRegs_1_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_1_4);
  assign multRegs_1_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_1_5);
  assign multRegs_1_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_1_6);
  assign multRegs_1_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_1_7);
  assign multRegs_1_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_1_8);
  assign multRegs_1_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_1_9);
  assign multRegs_1_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_1_10);
  assign multRegs_1_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_1_11);
  assign multRegs_1_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_1_12);
  assign multRegs_1_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_1_13);
  assign multRegs_1_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_1_14);
  assign multRegs_1_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_1_15);
  assign multRegs_2_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_2_0);
  assign multRegs_2_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_2_1);
  assign multRegs_2_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_2_2);
  assign multRegs_2_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_2_3);
  assign multRegs_2_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_2_4);
  assign multRegs_2_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_2_5);
  assign multRegs_2_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_2_6);
  assign multRegs_2_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_2_7);
  assign multRegs_2_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_2_8);
  assign multRegs_2_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_2_9);
  assign multRegs_2_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_2_10);
  assign multRegs_2_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_2_11);
  assign multRegs_2_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_2_12);
  assign multRegs_2_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_2_13);
  assign multRegs_2_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_2_14);
  assign multRegs_2_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_2_15);
  assign multRegs_3_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_3_0);
  assign multRegs_3_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_3_1);
  assign multRegs_3_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_3_2);
  assign multRegs_3_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_3_3);
  assign multRegs_3_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_3_4);
  assign multRegs_3_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_3_5);
  assign multRegs_3_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_3_6);
  assign multRegs_3_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_3_7);
  assign multRegs_3_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_3_8);
  assign multRegs_3_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_3_9);
  assign multRegs_3_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_3_10);
  assign multRegs_3_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_3_11);
  assign multRegs_3_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_3_12);
  assign multRegs_3_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_3_13);
  assign multRegs_3_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_3_14);
  assign multRegs_3_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_3_15);
  assign multRegs_4_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_4_0);
  assign multRegs_4_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_4_1);
  assign multRegs_4_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_4_2);
  assign multRegs_4_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_4_3);
  assign multRegs_4_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_4_4);
  assign multRegs_4_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_4_5);
  assign multRegs_4_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_4_6);
  assign multRegs_4_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_4_7);
  assign multRegs_4_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_4_8);
  assign multRegs_4_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_4_9);
  assign multRegs_4_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_4_10);
  assign multRegs_4_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_4_11);
  assign multRegs_4_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_4_12);
  assign multRegs_4_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_4_13);
  assign multRegs_4_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_4_14);
  assign multRegs_4_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_4_15);
  assign multRegs_5_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_5_0);
  assign multRegs_5_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_5_1);
  assign multRegs_5_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_5_2);
  assign multRegs_5_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_5_3);
  assign multRegs_5_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_5_4);
  assign multRegs_5_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_5_5);
  assign multRegs_5_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_5_6);
  assign multRegs_5_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_5_7);
  assign multRegs_5_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_5_8);
  assign multRegs_5_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_5_9);
  assign multRegs_5_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_5_10);
  assign multRegs_5_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_5_11);
  assign multRegs_5_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_5_12);
  assign multRegs_5_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_5_13);
  assign multRegs_5_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_5_14);
  assign multRegs_5_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_5_15);
  assign multRegs_6_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_6_0);
  assign multRegs_6_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_6_1);
  assign multRegs_6_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_6_2);
  assign multRegs_6_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_6_3);
  assign multRegs_6_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_6_4);
  assign multRegs_6_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_6_5);
  assign multRegs_6_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_6_6);
  assign multRegs_6_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_6_7);
  assign multRegs_6_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_6_8);
  assign multRegs_6_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_6_9);
  assign multRegs_6_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_6_10);
  assign multRegs_6_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_6_11);
  assign multRegs_6_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_6_12);
  assign multRegs_6_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_6_13);
  assign multRegs_6_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_6_14);
  assign multRegs_6_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_6_15);
  assign multRegs_7_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_7_0);
  assign multRegs_7_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_7_1);
  assign multRegs_7_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_7_2);
  assign multRegs_7_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_7_3);
  assign multRegs_7_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_7_4);
  assign multRegs_7_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_7_5);
  assign multRegs_7_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_7_6);
  assign multRegs_7_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_7_7);
  assign multRegs_7_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_7_8);
  assign multRegs_7_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_7_9);
  assign multRegs_7_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_7_10);
  assign multRegs_7_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_7_11);
  assign multRegs_7_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_7_12);
  assign multRegs_7_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_7_13);
  assign multRegs_7_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_7_14);
  assign multRegs_7_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_7_15);
  assign multRegs_8_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_8_0);
  assign multRegs_8_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_8_1);
  assign multRegs_8_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_8_2);
  assign multRegs_8_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_8_3);
  assign multRegs_8_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_8_4);
  assign multRegs_8_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_8_5);
  assign multRegs_8_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_8_6);
  assign multRegs_8_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_8_7);
  assign multRegs_8_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_8_8);
  assign multRegs_8_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_8_9);
  assign multRegs_8_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_8_10);
  assign multRegs_8_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_8_11);
  assign multRegs_8_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_8_12);
  assign multRegs_8_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_8_13);
  assign multRegs_8_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_8_14);
  assign multRegs_8_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_8_15);
  assign multRegs_9_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_9_0);
  assign multRegs_9_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_9_1);
  assign multRegs_9_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_9_2);
  assign multRegs_9_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_9_3);
  assign multRegs_9_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_9_4);
  assign multRegs_9_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_9_5);
  assign multRegs_9_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_9_6);
  assign multRegs_9_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_9_7);
  assign multRegs_9_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_9_8);
  assign multRegs_9_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_9_9);
  assign multRegs_9_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_9_10);
  assign multRegs_9_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_9_11);
  assign multRegs_9_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_9_12);
  assign multRegs_9_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_9_13);
  assign multRegs_9_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_9_14);
  assign multRegs_9_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_9_15);
  assign multRegs_10_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_10_0);
  assign multRegs_10_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_10_1);
  assign multRegs_10_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_10_2);
  assign multRegs_10_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_10_3);
  assign multRegs_10_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_10_4);
  assign multRegs_10_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_10_5);
  assign multRegs_10_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_10_6);
  assign multRegs_10_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_10_7);
  assign multRegs_10_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_10_8);
  assign multRegs_10_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_10_9);
  assign multRegs_10_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_10_10);
  assign multRegs_10_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_10_11);
  assign multRegs_10_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_10_12);
  assign multRegs_10_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_10_13);
  assign multRegs_10_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_10_14);
  assign multRegs_10_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_10_15);
  assign multRegs_11_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_11_0);
  assign multRegs_11_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_11_1);
  assign multRegs_11_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_11_2);
  assign multRegs_11_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_11_3);
  assign multRegs_11_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_11_4);
  assign multRegs_11_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_11_5);
  assign multRegs_11_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_11_6);
  assign multRegs_11_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_11_7);
  assign multRegs_11_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_11_8);
  assign multRegs_11_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_11_9);
  assign multRegs_11_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_11_10);
  assign multRegs_11_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_11_11);
  assign multRegs_11_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_11_12);
  assign multRegs_11_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_11_13);
  assign multRegs_11_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_11_14);
  assign multRegs_11_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_11_15);
  assign multRegs_12_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_12_0);
  assign multRegs_12_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_12_1);
  assign multRegs_12_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_12_2);
  assign multRegs_12_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_12_3);
  assign multRegs_12_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_12_4);
  assign multRegs_12_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_12_5);
  assign multRegs_12_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_12_6);
  assign multRegs_12_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_12_7);
  assign multRegs_12_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_12_8);
  assign multRegs_12_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_12_9);
  assign multRegs_12_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_12_10);
  assign multRegs_12_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_12_11);
  assign multRegs_12_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_12_12);
  assign multRegs_12_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_12_13);
  assign multRegs_12_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_12_14);
  assign multRegs_12_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_12_15);
  assign multRegs_13_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_13_0);
  assign multRegs_13_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_13_1);
  assign multRegs_13_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_13_2);
  assign multRegs_13_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_13_3);
  assign multRegs_13_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_13_4);
  assign multRegs_13_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_13_5);
  assign multRegs_13_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_13_6);
  assign multRegs_13_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_13_7);
  assign multRegs_13_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_13_8);
  assign multRegs_13_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_13_9);
  assign multRegs_13_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_13_10);
  assign multRegs_13_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_13_11);
  assign multRegs_13_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_13_12);
  assign multRegs_13_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_13_13);
  assign multRegs_13_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_13_14);
  assign multRegs_13_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_13_15);
  assign multRegs_14_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_14_0);
  assign multRegs_14_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_14_1);
  assign multRegs_14_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_14_2);
  assign multRegs_14_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_14_3);
  assign multRegs_14_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_14_4);
  assign multRegs_14_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_14_5);
  assign multRegs_14_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_14_6);
  assign multRegs_14_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_14_7);
  assign multRegs_14_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_14_8);
  assign multRegs_14_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_14_9);
  assign multRegs_14_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_14_10);
  assign multRegs_14_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_14_11);
  assign multRegs_14_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_14_12);
  assign multRegs_14_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_14_13);
  assign multRegs_14_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_14_14);
  assign multRegs_14_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_14_15);
  assign multRegs_15_0 = (io_inputDataIn_payload_0 * io_weightDataIn_payload_15_0);
  assign multRegs_15_1 = (io_inputDataIn_payload_1 * io_weightDataIn_payload_15_1);
  assign multRegs_15_2 = (io_inputDataIn_payload_2 * io_weightDataIn_payload_15_2);
  assign multRegs_15_3 = (io_inputDataIn_payload_3 * io_weightDataIn_payload_15_3);
  assign multRegs_15_4 = (io_inputDataIn_payload_4 * io_weightDataIn_payload_15_4);
  assign multRegs_15_5 = (io_inputDataIn_payload_5 * io_weightDataIn_payload_15_5);
  assign multRegs_15_6 = (io_inputDataIn_payload_6 * io_weightDataIn_payload_15_6);
  assign multRegs_15_7 = (io_inputDataIn_payload_7 * io_weightDataIn_payload_15_7);
  assign multRegs_15_8 = (io_inputDataIn_payload_8 * io_weightDataIn_payload_15_8);
  assign multRegs_15_9 = (io_inputDataIn_payload_9 * io_weightDataIn_payload_15_9);
  assign multRegs_15_10 = (io_inputDataIn_payload_10 * io_weightDataIn_payload_15_10);
  assign multRegs_15_11 = (io_inputDataIn_payload_11 * io_weightDataIn_payload_15_11);
  assign multRegs_15_12 = (io_inputDataIn_payload_12 * io_weightDataIn_payload_15_12);
  assign multRegs_15_13 = (io_inputDataIn_payload_13 * io_weightDataIn_payload_15_13);
  assign multRegs_15_14 = (io_inputDataIn_payload_14 * io_weightDataIn_payload_15_14);
  assign multRegs_15_15 = (io_inputDataIn_payload_15 * io_weightDataIn_payload_15_15);
  assign _zz_1 = ({1'b0,multRegs_0_0} + {1'b0,multRegs_0_8});
  assign _zz_2 = ({1'b0,multRegs_0_1} + {1'b0,multRegs_0_9});
  assign _zz_3 = ({1'b0,multRegs_0_2} + {1'b0,multRegs_0_10});
  assign _zz_4 = ({1'b0,multRegs_0_3} + {1'b0,multRegs_0_11});
  assign _zz_5 = ({1'b0,multRegs_0_4} + {1'b0,multRegs_0_12});
  assign _zz_6 = ({1'b0,multRegs_0_5} + {1'b0,multRegs_0_13});
  assign _zz_7 = ({1'b0,multRegs_0_6} + {1'b0,multRegs_0_14});
  assign _zz_8 = ({1'b0,multRegs_0_7} + {1'b0,multRegs_0_15});
  assign _zz_9 = ({1'b0,_zz_1_regNext} + {1'b0,_zz_5_regNext});
  assign _zz_10 = ({1'b0,_zz_2_regNext} + {1'b0,_zz_6_regNext});
  assign _zz_11 = ({1'b0,_zz_3_regNext} + {1'b0,_zz_7_regNext});
  assign _zz_12 = ({1'b0,_zz_4_regNext} + {1'b0,_zz_8_regNext});
  assign _zz_13 = ({1'b0,_zz_9_regNext} + {1'b0,_zz_11_regNext});
  assign _zz_14 = ({1'b0,_zz_10_regNext} + {1'b0,_zz_12_regNext});
  assign _zz_15 = ({1'b0,_zz_13_regNext} + {1'b0,_zz_14_regNext});
  assign adderTrees_0_result = _zz_15_regNext;
  assign _zz_16 = ({1'b0,multRegs_1_0} + {1'b0,multRegs_1_8});
  assign _zz_17 = ({1'b0,multRegs_1_1} + {1'b0,multRegs_1_9});
  assign _zz_18 = ({1'b0,multRegs_1_2} + {1'b0,multRegs_1_10});
  assign _zz_19 = ({1'b0,multRegs_1_3} + {1'b0,multRegs_1_11});
  assign _zz_20 = ({1'b0,multRegs_1_4} + {1'b0,multRegs_1_12});
  assign _zz_21 = ({1'b0,multRegs_1_5} + {1'b0,multRegs_1_13});
  assign _zz_22 = ({1'b0,multRegs_1_6} + {1'b0,multRegs_1_14});
  assign _zz_23 = ({1'b0,multRegs_1_7} + {1'b0,multRegs_1_15});
  assign _zz_24 = ({1'b0,_zz_16_regNext} + {1'b0,_zz_20_regNext});
  assign _zz_25 = ({1'b0,_zz_17_regNext} + {1'b0,_zz_21_regNext});
  assign _zz_26 = ({1'b0,_zz_18_regNext} + {1'b0,_zz_22_regNext});
  assign _zz_27 = ({1'b0,_zz_19_regNext} + {1'b0,_zz_23_regNext});
  assign _zz_28 = ({1'b0,_zz_24_regNext} + {1'b0,_zz_26_regNext});
  assign _zz_29 = ({1'b0,_zz_25_regNext} + {1'b0,_zz_27_regNext});
  assign _zz_30 = ({1'b0,_zz_28_regNext} + {1'b0,_zz_29_regNext});
  assign adderTrees_1_result = _zz_30_regNext;
  assign _zz_31 = ({1'b0,multRegs_2_0} + {1'b0,multRegs_2_8});
  assign _zz_32 = ({1'b0,multRegs_2_1} + {1'b0,multRegs_2_9});
  assign _zz_33 = ({1'b0,multRegs_2_2} + {1'b0,multRegs_2_10});
  assign _zz_34 = ({1'b0,multRegs_2_3} + {1'b0,multRegs_2_11});
  assign _zz_35 = ({1'b0,multRegs_2_4} + {1'b0,multRegs_2_12});
  assign _zz_36 = ({1'b0,multRegs_2_5} + {1'b0,multRegs_2_13});
  assign _zz_37 = ({1'b0,multRegs_2_6} + {1'b0,multRegs_2_14});
  assign _zz_38 = ({1'b0,multRegs_2_7} + {1'b0,multRegs_2_15});
  assign _zz_39 = ({1'b0,_zz_31_regNext} + {1'b0,_zz_35_regNext});
  assign _zz_40 = ({1'b0,_zz_32_regNext} + {1'b0,_zz_36_regNext});
  assign _zz_41 = ({1'b0,_zz_33_regNext} + {1'b0,_zz_37_regNext});
  assign _zz_42 = ({1'b0,_zz_34_regNext} + {1'b0,_zz_38_regNext});
  assign _zz_43 = ({1'b0,_zz_39_regNext} + {1'b0,_zz_41_regNext});
  assign _zz_44 = ({1'b0,_zz_40_regNext} + {1'b0,_zz_42_regNext});
  assign _zz_45 = ({1'b0,_zz_43_regNext} + {1'b0,_zz_44_regNext});
  assign adderTrees_2_result = _zz_45_regNext;
  assign _zz_46 = ({1'b0,multRegs_3_0} + {1'b0,multRegs_3_8});
  assign _zz_47 = ({1'b0,multRegs_3_1} + {1'b0,multRegs_3_9});
  assign _zz_48 = ({1'b0,multRegs_3_2} + {1'b0,multRegs_3_10});
  assign _zz_49 = ({1'b0,multRegs_3_3} + {1'b0,multRegs_3_11});
  assign _zz_50 = ({1'b0,multRegs_3_4} + {1'b0,multRegs_3_12});
  assign _zz_51 = ({1'b0,multRegs_3_5} + {1'b0,multRegs_3_13});
  assign _zz_52 = ({1'b0,multRegs_3_6} + {1'b0,multRegs_3_14});
  assign _zz_53 = ({1'b0,multRegs_3_7} + {1'b0,multRegs_3_15});
  assign _zz_54 = ({1'b0,_zz_46_regNext} + {1'b0,_zz_50_regNext});
  assign _zz_55 = ({1'b0,_zz_47_regNext} + {1'b0,_zz_51_regNext});
  assign _zz_56 = ({1'b0,_zz_48_regNext} + {1'b0,_zz_52_regNext});
  assign _zz_57 = ({1'b0,_zz_49_regNext} + {1'b0,_zz_53_regNext});
  assign _zz_58 = ({1'b0,_zz_54_regNext} + {1'b0,_zz_56_regNext});
  assign _zz_59 = ({1'b0,_zz_55_regNext} + {1'b0,_zz_57_regNext});
  assign _zz_60 = ({1'b0,_zz_58_regNext} + {1'b0,_zz_59_regNext});
  assign adderTrees_3_result = _zz_60_regNext;
  assign _zz_61 = ({1'b0,multRegs_4_0} + {1'b0,multRegs_4_8});
  assign _zz_62 = ({1'b0,multRegs_4_1} + {1'b0,multRegs_4_9});
  assign _zz_63 = ({1'b0,multRegs_4_2} + {1'b0,multRegs_4_10});
  assign _zz_64 = ({1'b0,multRegs_4_3} + {1'b0,multRegs_4_11});
  assign _zz_65 = ({1'b0,multRegs_4_4} + {1'b0,multRegs_4_12});
  assign _zz_66 = ({1'b0,multRegs_4_5} + {1'b0,multRegs_4_13});
  assign _zz_67 = ({1'b0,multRegs_4_6} + {1'b0,multRegs_4_14});
  assign _zz_68 = ({1'b0,multRegs_4_7} + {1'b0,multRegs_4_15});
  assign _zz_69 = ({1'b0,_zz_61_regNext} + {1'b0,_zz_65_regNext});
  assign _zz_70 = ({1'b0,_zz_62_regNext} + {1'b0,_zz_66_regNext});
  assign _zz_71 = ({1'b0,_zz_63_regNext} + {1'b0,_zz_67_regNext});
  assign _zz_72 = ({1'b0,_zz_64_regNext} + {1'b0,_zz_68_regNext});
  assign _zz_73 = ({1'b0,_zz_69_regNext} + {1'b0,_zz_71_regNext});
  assign _zz_74 = ({1'b0,_zz_70_regNext} + {1'b0,_zz_72_regNext});
  assign _zz_75 = ({1'b0,_zz_73_regNext} + {1'b0,_zz_74_regNext});
  assign adderTrees_4_result = _zz_75_regNext;
  assign _zz_76 = ({1'b0,multRegs_5_0} + {1'b0,multRegs_5_8});
  assign _zz_77 = ({1'b0,multRegs_5_1} + {1'b0,multRegs_5_9});
  assign _zz_78 = ({1'b0,multRegs_5_2} + {1'b0,multRegs_5_10});
  assign _zz_79 = ({1'b0,multRegs_5_3} + {1'b0,multRegs_5_11});
  assign _zz_80 = ({1'b0,multRegs_5_4} + {1'b0,multRegs_5_12});
  assign _zz_81 = ({1'b0,multRegs_5_5} + {1'b0,multRegs_5_13});
  assign _zz_82 = ({1'b0,multRegs_5_6} + {1'b0,multRegs_5_14});
  assign _zz_83 = ({1'b0,multRegs_5_7} + {1'b0,multRegs_5_15});
  assign _zz_84 = ({1'b0,_zz_76_regNext} + {1'b0,_zz_80_regNext});
  assign _zz_85 = ({1'b0,_zz_77_regNext} + {1'b0,_zz_81_regNext});
  assign _zz_86 = ({1'b0,_zz_78_regNext} + {1'b0,_zz_82_regNext});
  assign _zz_87 = ({1'b0,_zz_79_regNext} + {1'b0,_zz_83_regNext});
  assign _zz_88 = ({1'b0,_zz_84_regNext} + {1'b0,_zz_86_regNext});
  assign _zz_89 = ({1'b0,_zz_85_regNext} + {1'b0,_zz_87_regNext});
  assign _zz_90 = ({1'b0,_zz_88_regNext} + {1'b0,_zz_89_regNext});
  assign adderTrees_5_result = _zz_90_regNext;
  assign _zz_91 = ({1'b0,multRegs_6_0} + {1'b0,multRegs_6_8});
  assign _zz_92 = ({1'b0,multRegs_6_1} + {1'b0,multRegs_6_9});
  assign _zz_93 = ({1'b0,multRegs_6_2} + {1'b0,multRegs_6_10});
  assign _zz_94 = ({1'b0,multRegs_6_3} + {1'b0,multRegs_6_11});
  assign _zz_95 = ({1'b0,multRegs_6_4} + {1'b0,multRegs_6_12});
  assign _zz_96 = ({1'b0,multRegs_6_5} + {1'b0,multRegs_6_13});
  assign _zz_97 = ({1'b0,multRegs_6_6} + {1'b0,multRegs_6_14});
  assign _zz_98 = ({1'b0,multRegs_6_7} + {1'b0,multRegs_6_15});
  assign _zz_99 = ({1'b0,_zz_91_regNext} + {1'b0,_zz_95_regNext});
  assign _zz_100 = ({1'b0,_zz_92_regNext} + {1'b0,_zz_96_regNext});
  assign _zz_101 = ({1'b0,_zz_93_regNext} + {1'b0,_zz_97_regNext});
  assign _zz_102 = ({1'b0,_zz_94_regNext} + {1'b0,_zz_98_regNext});
  assign _zz_103 = ({1'b0,_zz_99_regNext} + {1'b0,_zz_101_regNext});
  assign _zz_104 = ({1'b0,_zz_100_regNext} + {1'b0,_zz_102_regNext});
  assign _zz_105 = ({1'b0,_zz_103_regNext} + {1'b0,_zz_104_regNext});
  assign adderTrees_6_result = _zz_105_regNext;
  assign _zz_106 = ({1'b0,multRegs_7_0} + {1'b0,multRegs_7_8});
  assign _zz_107 = ({1'b0,multRegs_7_1} + {1'b0,multRegs_7_9});
  assign _zz_108 = ({1'b0,multRegs_7_2} + {1'b0,multRegs_7_10});
  assign _zz_109 = ({1'b0,multRegs_7_3} + {1'b0,multRegs_7_11});
  assign _zz_110 = ({1'b0,multRegs_7_4} + {1'b0,multRegs_7_12});
  assign _zz_111 = ({1'b0,multRegs_7_5} + {1'b0,multRegs_7_13});
  assign _zz_112 = ({1'b0,multRegs_7_6} + {1'b0,multRegs_7_14});
  assign _zz_113 = ({1'b0,multRegs_7_7} + {1'b0,multRegs_7_15});
  assign _zz_114 = ({1'b0,_zz_106_regNext} + {1'b0,_zz_110_regNext});
  assign _zz_115 = ({1'b0,_zz_107_regNext} + {1'b0,_zz_111_regNext});
  assign _zz_116 = ({1'b0,_zz_108_regNext} + {1'b0,_zz_112_regNext});
  assign _zz_117 = ({1'b0,_zz_109_regNext} + {1'b0,_zz_113_regNext});
  assign _zz_118 = ({1'b0,_zz_114_regNext} + {1'b0,_zz_116_regNext});
  assign _zz_119 = ({1'b0,_zz_115_regNext} + {1'b0,_zz_117_regNext});
  assign _zz_120 = ({1'b0,_zz_118_regNext} + {1'b0,_zz_119_regNext});
  assign adderTrees_7_result = _zz_120_regNext;
  assign _zz_121 = ({1'b0,multRegs_8_0} + {1'b0,multRegs_8_8});
  assign _zz_122 = ({1'b0,multRegs_8_1} + {1'b0,multRegs_8_9});
  assign _zz_123 = ({1'b0,multRegs_8_2} + {1'b0,multRegs_8_10});
  assign _zz_124 = ({1'b0,multRegs_8_3} + {1'b0,multRegs_8_11});
  assign _zz_125 = ({1'b0,multRegs_8_4} + {1'b0,multRegs_8_12});
  assign _zz_126 = ({1'b0,multRegs_8_5} + {1'b0,multRegs_8_13});
  assign _zz_127 = ({1'b0,multRegs_8_6} + {1'b0,multRegs_8_14});
  assign _zz_128 = ({1'b0,multRegs_8_7} + {1'b0,multRegs_8_15});
  assign _zz_129 = ({1'b0,_zz_121_regNext} + {1'b0,_zz_125_regNext});
  assign _zz_130 = ({1'b0,_zz_122_regNext} + {1'b0,_zz_126_regNext});
  assign _zz_131 = ({1'b0,_zz_123_regNext} + {1'b0,_zz_127_regNext});
  assign _zz_132 = ({1'b0,_zz_124_regNext} + {1'b0,_zz_128_regNext});
  assign _zz_133 = ({1'b0,_zz_129_regNext} + {1'b0,_zz_131_regNext});
  assign _zz_134 = ({1'b0,_zz_130_regNext} + {1'b0,_zz_132_regNext});
  assign _zz_135 = ({1'b0,_zz_133_regNext} + {1'b0,_zz_134_regNext});
  assign adderTrees_8_result = _zz_135_regNext;
  assign _zz_136 = ({1'b0,multRegs_9_0} + {1'b0,multRegs_9_8});
  assign _zz_137 = ({1'b0,multRegs_9_1} + {1'b0,multRegs_9_9});
  assign _zz_138 = ({1'b0,multRegs_9_2} + {1'b0,multRegs_9_10});
  assign _zz_139 = ({1'b0,multRegs_9_3} + {1'b0,multRegs_9_11});
  assign _zz_140 = ({1'b0,multRegs_9_4} + {1'b0,multRegs_9_12});
  assign _zz_141 = ({1'b0,multRegs_9_5} + {1'b0,multRegs_9_13});
  assign _zz_142 = ({1'b0,multRegs_9_6} + {1'b0,multRegs_9_14});
  assign _zz_143 = ({1'b0,multRegs_9_7} + {1'b0,multRegs_9_15});
  assign _zz_144 = ({1'b0,_zz_136_regNext} + {1'b0,_zz_140_regNext});
  assign _zz_145 = ({1'b0,_zz_137_regNext} + {1'b0,_zz_141_regNext});
  assign _zz_146 = ({1'b0,_zz_138_regNext} + {1'b0,_zz_142_regNext});
  assign _zz_147 = ({1'b0,_zz_139_regNext} + {1'b0,_zz_143_regNext});
  assign _zz_148 = ({1'b0,_zz_144_regNext} + {1'b0,_zz_146_regNext});
  assign _zz_149 = ({1'b0,_zz_145_regNext} + {1'b0,_zz_147_regNext});
  assign _zz_150 = ({1'b0,_zz_148_regNext} + {1'b0,_zz_149_regNext});
  assign adderTrees_9_result = _zz_150_regNext;
  assign _zz_151 = ({1'b0,multRegs_10_0} + {1'b0,multRegs_10_8});
  assign _zz_152 = ({1'b0,multRegs_10_1} + {1'b0,multRegs_10_9});
  assign _zz_153 = ({1'b0,multRegs_10_2} + {1'b0,multRegs_10_10});
  assign _zz_154 = ({1'b0,multRegs_10_3} + {1'b0,multRegs_10_11});
  assign _zz_155 = ({1'b0,multRegs_10_4} + {1'b0,multRegs_10_12});
  assign _zz_156 = ({1'b0,multRegs_10_5} + {1'b0,multRegs_10_13});
  assign _zz_157 = ({1'b0,multRegs_10_6} + {1'b0,multRegs_10_14});
  assign _zz_158 = ({1'b0,multRegs_10_7} + {1'b0,multRegs_10_15});
  assign _zz_159 = ({1'b0,_zz_151_regNext} + {1'b0,_zz_155_regNext});
  assign _zz_160 = ({1'b0,_zz_152_regNext} + {1'b0,_zz_156_regNext});
  assign _zz_161 = ({1'b0,_zz_153_regNext} + {1'b0,_zz_157_regNext});
  assign _zz_162 = ({1'b0,_zz_154_regNext} + {1'b0,_zz_158_regNext});
  assign _zz_163 = ({1'b0,_zz_159_regNext} + {1'b0,_zz_161_regNext});
  assign _zz_164 = ({1'b0,_zz_160_regNext} + {1'b0,_zz_162_regNext});
  assign _zz_165 = ({1'b0,_zz_163_regNext} + {1'b0,_zz_164_regNext});
  assign adderTrees_10_result = _zz_165_regNext;
  assign _zz_166 = ({1'b0,multRegs_11_0} + {1'b0,multRegs_11_8});
  assign _zz_167 = ({1'b0,multRegs_11_1} + {1'b0,multRegs_11_9});
  assign _zz_168 = ({1'b0,multRegs_11_2} + {1'b0,multRegs_11_10});
  assign _zz_169 = ({1'b0,multRegs_11_3} + {1'b0,multRegs_11_11});
  assign _zz_170 = ({1'b0,multRegs_11_4} + {1'b0,multRegs_11_12});
  assign _zz_171 = ({1'b0,multRegs_11_5} + {1'b0,multRegs_11_13});
  assign _zz_172 = ({1'b0,multRegs_11_6} + {1'b0,multRegs_11_14});
  assign _zz_173 = ({1'b0,multRegs_11_7} + {1'b0,multRegs_11_15});
  assign _zz_174 = ({1'b0,_zz_166_regNext} + {1'b0,_zz_170_regNext});
  assign _zz_175 = ({1'b0,_zz_167_regNext} + {1'b0,_zz_171_regNext});
  assign _zz_176 = ({1'b0,_zz_168_regNext} + {1'b0,_zz_172_regNext});
  assign _zz_177 = ({1'b0,_zz_169_regNext} + {1'b0,_zz_173_regNext});
  assign _zz_178 = ({1'b0,_zz_174_regNext} + {1'b0,_zz_176_regNext});
  assign _zz_179 = ({1'b0,_zz_175_regNext} + {1'b0,_zz_177_regNext});
  assign _zz_180 = ({1'b0,_zz_178_regNext} + {1'b0,_zz_179_regNext});
  assign adderTrees_11_result = _zz_180_regNext;
  assign _zz_181 = ({1'b0,multRegs_12_0} + {1'b0,multRegs_12_8});
  assign _zz_182 = ({1'b0,multRegs_12_1} + {1'b0,multRegs_12_9});
  assign _zz_183 = ({1'b0,multRegs_12_2} + {1'b0,multRegs_12_10});
  assign _zz_184 = ({1'b0,multRegs_12_3} + {1'b0,multRegs_12_11});
  assign _zz_185 = ({1'b0,multRegs_12_4} + {1'b0,multRegs_12_12});
  assign _zz_186 = ({1'b0,multRegs_12_5} + {1'b0,multRegs_12_13});
  assign _zz_187 = ({1'b0,multRegs_12_6} + {1'b0,multRegs_12_14});
  assign _zz_188 = ({1'b0,multRegs_12_7} + {1'b0,multRegs_12_15});
  assign _zz_189 = ({1'b0,_zz_181_regNext} + {1'b0,_zz_185_regNext});
  assign _zz_190 = ({1'b0,_zz_182_regNext} + {1'b0,_zz_186_regNext});
  assign _zz_191 = ({1'b0,_zz_183_regNext} + {1'b0,_zz_187_regNext});
  assign _zz_192 = ({1'b0,_zz_184_regNext} + {1'b0,_zz_188_regNext});
  assign _zz_193 = ({1'b0,_zz_189_regNext} + {1'b0,_zz_191_regNext});
  assign _zz_194 = ({1'b0,_zz_190_regNext} + {1'b0,_zz_192_regNext});
  assign _zz_195 = ({1'b0,_zz_193_regNext} + {1'b0,_zz_194_regNext});
  assign adderTrees_12_result = _zz_195_regNext;
  assign _zz_196 = ({1'b0,multRegs_13_0} + {1'b0,multRegs_13_8});
  assign _zz_197 = ({1'b0,multRegs_13_1} + {1'b0,multRegs_13_9});
  assign _zz_198 = ({1'b0,multRegs_13_2} + {1'b0,multRegs_13_10});
  assign _zz_199 = ({1'b0,multRegs_13_3} + {1'b0,multRegs_13_11});
  assign _zz_200 = ({1'b0,multRegs_13_4} + {1'b0,multRegs_13_12});
  assign _zz_201 = ({1'b0,multRegs_13_5} + {1'b0,multRegs_13_13});
  assign _zz_202 = ({1'b0,multRegs_13_6} + {1'b0,multRegs_13_14});
  assign _zz_203 = ({1'b0,multRegs_13_7} + {1'b0,multRegs_13_15});
  assign _zz_204 = ({1'b0,_zz_196_regNext} + {1'b0,_zz_200_regNext});
  assign _zz_205 = ({1'b0,_zz_197_regNext} + {1'b0,_zz_201_regNext});
  assign _zz_206 = ({1'b0,_zz_198_regNext} + {1'b0,_zz_202_regNext});
  assign _zz_207 = ({1'b0,_zz_199_regNext} + {1'b0,_zz_203_regNext});
  assign _zz_208 = ({1'b0,_zz_204_regNext} + {1'b0,_zz_206_regNext});
  assign _zz_209 = ({1'b0,_zz_205_regNext} + {1'b0,_zz_207_regNext});
  assign _zz_210 = ({1'b0,_zz_208_regNext} + {1'b0,_zz_209_regNext});
  assign adderTrees_13_result = _zz_210_regNext;
  assign _zz_211 = ({1'b0,multRegs_14_0} + {1'b0,multRegs_14_8});
  assign _zz_212 = ({1'b0,multRegs_14_1} + {1'b0,multRegs_14_9});
  assign _zz_213 = ({1'b0,multRegs_14_2} + {1'b0,multRegs_14_10});
  assign _zz_214 = ({1'b0,multRegs_14_3} + {1'b0,multRegs_14_11});
  assign _zz_215 = ({1'b0,multRegs_14_4} + {1'b0,multRegs_14_12});
  assign _zz_216 = ({1'b0,multRegs_14_5} + {1'b0,multRegs_14_13});
  assign _zz_217 = ({1'b0,multRegs_14_6} + {1'b0,multRegs_14_14});
  assign _zz_218 = ({1'b0,multRegs_14_7} + {1'b0,multRegs_14_15});
  assign _zz_219 = ({1'b0,_zz_211_regNext} + {1'b0,_zz_215_regNext});
  assign _zz_220 = ({1'b0,_zz_212_regNext} + {1'b0,_zz_216_regNext});
  assign _zz_221 = ({1'b0,_zz_213_regNext} + {1'b0,_zz_217_regNext});
  assign _zz_222 = ({1'b0,_zz_214_regNext} + {1'b0,_zz_218_regNext});
  assign _zz_223 = ({1'b0,_zz_219_regNext} + {1'b0,_zz_221_regNext});
  assign _zz_224 = ({1'b0,_zz_220_regNext} + {1'b0,_zz_222_regNext});
  assign _zz_225 = ({1'b0,_zz_223_regNext} + {1'b0,_zz_224_regNext});
  assign adderTrees_14_result = _zz_225_regNext;
  assign _zz_226 = ({1'b0,multRegs_15_0} + {1'b0,multRegs_15_8});
  assign _zz_227 = ({1'b0,multRegs_15_1} + {1'b0,multRegs_15_9});
  assign _zz_228 = ({1'b0,multRegs_15_2} + {1'b0,multRegs_15_10});
  assign _zz_229 = ({1'b0,multRegs_15_3} + {1'b0,multRegs_15_11});
  assign _zz_230 = ({1'b0,multRegs_15_4} + {1'b0,multRegs_15_12});
  assign _zz_231 = ({1'b0,multRegs_15_5} + {1'b0,multRegs_15_13});
  assign _zz_232 = ({1'b0,multRegs_15_6} + {1'b0,multRegs_15_14});
  assign _zz_233 = ({1'b0,multRegs_15_7} + {1'b0,multRegs_15_15});
  assign _zz_234 = ({1'b0,_zz_226_regNext} + {1'b0,_zz_230_regNext});
  assign _zz_235 = ({1'b0,_zz_227_regNext} + {1'b0,_zz_231_regNext});
  assign _zz_236 = ({1'b0,_zz_228_regNext} + {1'b0,_zz_232_regNext});
  assign _zz_237 = ({1'b0,_zz_229_regNext} + {1'b0,_zz_233_regNext});
  assign _zz_238 = ({1'b0,_zz_234_regNext} + {1'b0,_zz_236_regNext});
  assign _zz_239 = ({1'b0,_zz_235_regNext} + {1'b0,_zz_237_regNext});
  assign _zz_240 = ({1'b0,_zz_238_regNext} + {1'b0,_zz_239_regNext});
  assign adderTrees_15_result = _zz_240_regNext;
  assign io_inputDataIn_ready = io_calc2write_1_ready;
  assign io_weightDataIn_ready = io_calc2write_1_ready;
  always @ (*) begin
    validCounter_willIncrement = 1'b0;
    if(((io_inputDataIn_valid && io_inputDataIn_ready) && (io_weightDataIn_valid && io_weightDataIn_ready)))begin
      validCounter_willIncrement = 1'b1;
    end
  end

  assign validCounter_willClear = 1'b0;
  assign validCounter_willOverflowIfInc = (validCounter_value == 2'b11);
  assign validCounter_willOverflow = (validCounter_willOverflowIfInc && validCounter_willIncrement);
  always @ (*) begin
    validCounter_valueNext = (validCounter_value + _zz_242);
    if(validCounter_willClear)begin
      validCounter_valueNext = 2'b00;
    end
  end

  assign io_calc2write_1_payload_0 = accRegs_0[7:0];
  assign io_calc2write_1_payload_1 = accRegs_1[7:0];
  assign io_calc2write_1_payload_2 = accRegs_2[7:0];
  assign io_calc2write_1_payload_3 = accRegs_3[7:0];
  assign io_calc2write_1_payload_4 = accRegs_4[7:0];
  assign io_calc2write_1_payload_5 = accRegs_5[7:0];
  assign io_calc2write_1_payload_6 = accRegs_6[7:0];
  assign io_calc2write_1_payload_7 = accRegs_7[7:0];
  assign io_calc2write_1_payload_8 = accRegs_8[7:0];
  assign io_calc2write_1_payload_9 = accRegs_9[7:0];
  assign io_calc2write_1_payload_10 = accRegs_10[7:0];
  assign io_calc2write_1_payload_11 = accRegs_11[7:0];
  assign io_calc2write_1_payload_12 = accRegs_12[7:0];
  assign io_calc2write_1_payload_13 = accRegs_13[7:0];
  assign io_calc2write_1_payload_14 = accRegs_14[7:0];
  assign io_calc2write_1_payload_15 = accRegs_15[7:0];
  assign io_calc2write_1_valid = validCounter_willOverflow_delay_5;
  always @ (posedge clk) begin
    _zz_1_regNext <= _zz_1;
    _zz_2_regNext <= _zz_2;
    _zz_3_regNext <= _zz_3;
    _zz_4_regNext <= _zz_4;
    _zz_5_regNext <= _zz_5;
    _zz_6_regNext <= _zz_6;
    _zz_7_regNext <= _zz_7;
    _zz_8_regNext <= _zz_8;
    _zz_9_regNext <= _zz_9;
    _zz_10_regNext <= _zz_10;
    _zz_11_regNext <= _zz_11;
    _zz_12_regNext <= _zz_12;
    _zz_13_regNext <= _zz_13;
    _zz_14_regNext <= _zz_14;
    _zz_15_regNext <= _zz_15;
    _zz_16_regNext <= _zz_16;
    _zz_17_regNext <= _zz_17;
    _zz_18_regNext <= _zz_18;
    _zz_19_regNext <= _zz_19;
    _zz_20_regNext <= _zz_20;
    _zz_21_regNext <= _zz_21;
    _zz_22_regNext <= _zz_22;
    _zz_23_regNext <= _zz_23;
    _zz_24_regNext <= _zz_24;
    _zz_25_regNext <= _zz_25;
    _zz_26_regNext <= _zz_26;
    _zz_27_regNext <= _zz_27;
    _zz_28_regNext <= _zz_28;
    _zz_29_regNext <= _zz_29;
    _zz_30_regNext <= _zz_30;
    _zz_31_regNext <= _zz_31;
    _zz_32_regNext <= _zz_32;
    _zz_33_regNext <= _zz_33;
    _zz_34_regNext <= _zz_34;
    _zz_35_regNext <= _zz_35;
    _zz_36_regNext <= _zz_36;
    _zz_37_regNext <= _zz_37;
    _zz_38_regNext <= _zz_38;
    _zz_39_regNext <= _zz_39;
    _zz_40_regNext <= _zz_40;
    _zz_41_regNext <= _zz_41;
    _zz_42_regNext <= _zz_42;
    _zz_43_regNext <= _zz_43;
    _zz_44_regNext <= _zz_44;
    _zz_45_regNext <= _zz_45;
    _zz_46_regNext <= _zz_46;
    _zz_47_regNext <= _zz_47;
    _zz_48_regNext <= _zz_48;
    _zz_49_regNext <= _zz_49;
    _zz_50_regNext <= _zz_50;
    _zz_51_regNext <= _zz_51;
    _zz_52_regNext <= _zz_52;
    _zz_53_regNext <= _zz_53;
    _zz_54_regNext <= _zz_54;
    _zz_55_regNext <= _zz_55;
    _zz_56_regNext <= _zz_56;
    _zz_57_regNext <= _zz_57;
    _zz_58_regNext <= _zz_58;
    _zz_59_regNext <= _zz_59;
    _zz_60_regNext <= _zz_60;
    _zz_61_regNext <= _zz_61;
    _zz_62_regNext <= _zz_62;
    _zz_63_regNext <= _zz_63;
    _zz_64_regNext <= _zz_64;
    _zz_65_regNext <= _zz_65;
    _zz_66_regNext <= _zz_66;
    _zz_67_regNext <= _zz_67;
    _zz_68_regNext <= _zz_68;
    _zz_69_regNext <= _zz_69;
    _zz_70_regNext <= _zz_70;
    _zz_71_regNext <= _zz_71;
    _zz_72_regNext <= _zz_72;
    _zz_73_regNext <= _zz_73;
    _zz_74_regNext <= _zz_74;
    _zz_75_regNext <= _zz_75;
    _zz_76_regNext <= _zz_76;
    _zz_77_regNext <= _zz_77;
    _zz_78_regNext <= _zz_78;
    _zz_79_regNext <= _zz_79;
    _zz_80_regNext <= _zz_80;
    _zz_81_regNext <= _zz_81;
    _zz_82_regNext <= _zz_82;
    _zz_83_regNext <= _zz_83;
    _zz_84_regNext <= _zz_84;
    _zz_85_regNext <= _zz_85;
    _zz_86_regNext <= _zz_86;
    _zz_87_regNext <= _zz_87;
    _zz_88_regNext <= _zz_88;
    _zz_89_regNext <= _zz_89;
    _zz_90_regNext <= _zz_90;
    _zz_91_regNext <= _zz_91;
    _zz_92_regNext <= _zz_92;
    _zz_93_regNext <= _zz_93;
    _zz_94_regNext <= _zz_94;
    _zz_95_regNext <= _zz_95;
    _zz_96_regNext <= _zz_96;
    _zz_97_regNext <= _zz_97;
    _zz_98_regNext <= _zz_98;
    _zz_99_regNext <= _zz_99;
    _zz_100_regNext <= _zz_100;
    _zz_101_regNext <= _zz_101;
    _zz_102_regNext <= _zz_102;
    _zz_103_regNext <= _zz_103;
    _zz_104_regNext <= _zz_104;
    _zz_105_regNext <= _zz_105;
    _zz_106_regNext <= _zz_106;
    _zz_107_regNext <= _zz_107;
    _zz_108_regNext <= _zz_108;
    _zz_109_regNext <= _zz_109;
    _zz_110_regNext <= _zz_110;
    _zz_111_regNext <= _zz_111;
    _zz_112_regNext <= _zz_112;
    _zz_113_regNext <= _zz_113;
    _zz_114_regNext <= _zz_114;
    _zz_115_regNext <= _zz_115;
    _zz_116_regNext <= _zz_116;
    _zz_117_regNext <= _zz_117;
    _zz_118_regNext <= _zz_118;
    _zz_119_regNext <= _zz_119;
    _zz_120_regNext <= _zz_120;
    _zz_121_regNext <= _zz_121;
    _zz_122_regNext <= _zz_122;
    _zz_123_regNext <= _zz_123;
    _zz_124_regNext <= _zz_124;
    _zz_125_regNext <= _zz_125;
    _zz_126_regNext <= _zz_126;
    _zz_127_regNext <= _zz_127;
    _zz_128_regNext <= _zz_128;
    _zz_129_regNext <= _zz_129;
    _zz_130_regNext <= _zz_130;
    _zz_131_regNext <= _zz_131;
    _zz_132_regNext <= _zz_132;
    _zz_133_regNext <= _zz_133;
    _zz_134_regNext <= _zz_134;
    _zz_135_regNext <= _zz_135;
    _zz_136_regNext <= _zz_136;
    _zz_137_regNext <= _zz_137;
    _zz_138_regNext <= _zz_138;
    _zz_139_regNext <= _zz_139;
    _zz_140_regNext <= _zz_140;
    _zz_141_regNext <= _zz_141;
    _zz_142_regNext <= _zz_142;
    _zz_143_regNext <= _zz_143;
    _zz_144_regNext <= _zz_144;
    _zz_145_regNext <= _zz_145;
    _zz_146_regNext <= _zz_146;
    _zz_147_regNext <= _zz_147;
    _zz_148_regNext <= _zz_148;
    _zz_149_regNext <= _zz_149;
    _zz_150_regNext <= _zz_150;
    _zz_151_regNext <= _zz_151;
    _zz_152_regNext <= _zz_152;
    _zz_153_regNext <= _zz_153;
    _zz_154_regNext <= _zz_154;
    _zz_155_regNext <= _zz_155;
    _zz_156_regNext <= _zz_156;
    _zz_157_regNext <= _zz_157;
    _zz_158_regNext <= _zz_158;
    _zz_159_regNext <= _zz_159;
    _zz_160_regNext <= _zz_160;
    _zz_161_regNext <= _zz_161;
    _zz_162_regNext <= _zz_162;
    _zz_163_regNext <= _zz_163;
    _zz_164_regNext <= _zz_164;
    _zz_165_regNext <= _zz_165;
    _zz_166_regNext <= _zz_166;
    _zz_167_regNext <= _zz_167;
    _zz_168_regNext <= _zz_168;
    _zz_169_regNext <= _zz_169;
    _zz_170_regNext <= _zz_170;
    _zz_171_regNext <= _zz_171;
    _zz_172_regNext <= _zz_172;
    _zz_173_regNext <= _zz_173;
    _zz_174_regNext <= _zz_174;
    _zz_175_regNext <= _zz_175;
    _zz_176_regNext <= _zz_176;
    _zz_177_regNext <= _zz_177;
    _zz_178_regNext <= _zz_178;
    _zz_179_regNext <= _zz_179;
    _zz_180_regNext <= _zz_180;
    _zz_181_regNext <= _zz_181;
    _zz_182_regNext <= _zz_182;
    _zz_183_regNext <= _zz_183;
    _zz_184_regNext <= _zz_184;
    _zz_185_regNext <= _zz_185;
    _zz_186_regNext <= _zz_186;
    _zz_187_regNext <= _zz_187;
    _zz_188_regNext <= _zz_188;
    _zz_189_regNext <= _zz_189;
    _zz_190_regNext <= _zz_190;
    _zz_191_regNext <= _zz_191;
    _zz_192_regNext <= _zz_192;
    _zz_193_regNext <= _zz_193;
    _zz_194_regNext <= _zz_194;
    _zz_195_regNext <= _zz_195;
    _zz_196_regNext <= _zz_196;
    _zz_197_regNext <= _zz_197;
    _zz_198_regNext <= _zz_198;
    _zz_199_regNext <= _zz_199;
    _zz_200_regNext <= _zz_200;
    _zz_201_regNext <= _zz_201;
    _zz_202_regNext <= _zz_202;
    _zz_203_regNext <= _zz_203;
    _zz_204_regNext <= _zz_204;
    _zz_205_regNext <= _zz_205;
    _zz_206_regNext <= _zz_206;
    _zz_207_regNext <= _zz_207;
    _zz_208_regNext <= _zz_208;
    _zz_209_regNext <= _zz_209;
    _zz_210_regNext <= _zz_210;
    _zz_211_regNext <= _zz_211;
    _zz_212_regNext <= _zz_212;
    _zz_213_regNext <= _zz_213;
    _zz_214_regNext <= _zz_214;
    _zz_215_regNext <= _zz_215;
    _zz_216_regNext <= _zz_216;
    _zz_217_regNext <= _zz_217;
    _zz_218_regNext <= _zz_218;
    _zz_219_regNext <= _zz_219;
    _zz_220_regNext <= _zz_220;
    _zz_221_regNext <= _zz_221;
    _zz_222_regNext <= _zz_222;
    _zz_223_regNext <= _zz_223;
    _zz_224_regNext <= _zz_224;
    _zz_225_regNext <= _zz_225;
    _zz_226_regNext <= _zz_226;
    _zz_227_regNext <= _zz_227;
    _zz_228_regNext <= _zz_228;
    _zz_229_regNext <= _zz_229;
    _zz_230_regNext <= _zz_230;
    _zz_231_regNext <= _zz_231;
    _zz_232_regNext <= _zz_232;
    _zz_233_regNext <= _zz_233;
    _zz_234_regNext <= _zz_234;
    _zz_235_regNext <= _zz_235;
    _zz_236_regNext <= _zz_236;
    _zz_237_regNext <= _zz_237;
    _zz_238_regNext <= _zz_238;
    _zz_239_regNext <= _zz_239;
    _zz_240_regNext <= _zz_240;
    if(validCounter_willOverflow)begin
      accRegs_0 <= {2'd0, adderTrees_0_result};
      accRegs_1 <= {2'd0, adderTrees_1_result};
      accRegs_2 <= {2'd0, adderTrees_2_result};
      accRegs_3 <= {2'd0, adderTrees_3_result};
      accRegs_4 <= {2'd0, adderTrees_4_result};
      accRegs_5 <= {2'd0, adderTrees_5_result};
      accRegs_6 <= {2'd0, adderTrees_6_result};
      accRegs_7 <= {2'd0, adderTrees_7_result};
      accRegs_8 <= {2'd0, adderTrees_8_result};
      accRegs_9 <= {2'd0, adderTrees_9_result};
      accRegs_10 <= {2'd0, adderTrees_10_result};
      accRegs_11 <= {2'd0, adderTrees_11_result};
      accRegs_12 <= {2'd0, adderTrees_12_result};
      accRegs_13 <= {2'd0, adderTrees_13_result};
      accRegs_14 <= {2'd0, adderTrees_14_result};
      accRegs_15 <= {2'd0, adderTrees_15_result};
    end else begin
      accRegs_0 <= (accRegs_0 + _zz_243);
      accRegs_1 <= (accRegs_1 + _zz_244);
      accRegs_2 <= (accRegs_2 + _zz_245);
      accRegs_3 <= (accRegs_3 + _zz_246);
      accRegs_4 <= (accRegs_4 + _zz_247);
      accRegs_5 <= (accRegs_5 + _zz_248);
      accRegs_6 <= (accRegs_6 + _zz_249);
      accRegs_7 <= (accRegs_7 + _zz_250);
      accRegs_8 <= (accRegs_8 + _zz_251);
      accRegs_9 <= (accRegs_9 + _zz_252);
      accRegs_10 <= (accRegs_10 + _zz_253);
      accRegs_11 <= (accRegs_11 + _zz_254);
      accRegs_12 <= (accRegs_12 + _zz_255);
      accRegs_13 <= (accRegs_13 + _zz_256);
      accRegs_14 <= (accRegs_14 + _zz_257);
      accRegs_15 <= (accRegs_15 + _zz_258);
    end
    validCounter_willOverflow_delay_1 <= validCounter_willOverflow;
    validCounter_willOverflow_delay_2 <= validCounter_willOverflow_delay_1;
    validCounter_willOverflow_delay_3 <= validCounter_willOverflow_delay_2;
    validCounter_willOverflow_delay_4 <= validCounter_willOverflow_delay_3;
    validCounter_willOverflow_delay_5 <= validCounter_willOverflow_delay_4;
  end

  always @ (posedge clk or posedge reset) begin
    if (reset) begin
      validCounter_value <= 2'b00;
    end else begin
      validCounter_value <= validCounter_valueNext;
    end
  end


endmodule
